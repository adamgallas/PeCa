// Generator : SpinalHDL v1.6.4    git head : 598c18959149eb18e5eee5b0aa3eef01ecaa41a1
// Component : PeCa

`timescale 1ns/1ps 

module PeCa (
  input      [7:0]    numberOfInputFrames,
  input      [7:0]    numberOfOutputFrames,
  input      [8:0]    width,
  input      [8:0]    height,
  input      [7:0]    inputZeroPoint,
  input      [7:0]    outputZeroPoint,
  input      [15:0]   scaleBase,
  input      [5:0]    scaleExpr,
  input               enablePooling,
  input               inputs_valid,
  output              inputs_ready,
  input      [127:0]  inputs_payload,
  input               weights_valid,
  output              weights_ready,
  input      [127:0]  weights_payload,
  input               funcTable_valid,
  output              funcTable_ready,
  input      [127:0]  funcTable_payload,
  output              outputs_valid,
  input               outputs_ready,
  output     [127:0]  outputs_payload,
  input               clk,
  input               reset
);

  wire       [0:0]    streamDemux_3_io_select;
  wire       [0:0]    streamMux_1_io_select;
  wire                weightFifo_0_push_ready;
  wire                weightFifo_0_pop_valid;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_0_pop_payload_1_2_2_15;
  wire                weightFifo_1_push_ready;
  wire                weightFifo_1_pop_valid;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_1_pop_payload_1_2_2_15;
  wire                weightFifo_2_push_ready;
  wire                weightFifo_2_pop_valid;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_2_pop_payload_1_2_2_15;
  wire                weightFifo_3_push_ready;
  wire                weightFifo_3_pop_valid;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_3_pop_payload_1_2_2_15;
  wire                weightFifo_4_push_ready;
  wire                weightFifo_4_pop_valid;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_4_pop_payload_1_2_2_15;
  wire                weightFifo_5_push_ready;
  wire                weightFifo_5_pop_valid;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_5_pop_payload_1_2_2_15;
  wire                weightFifo_6_push_ready;
  wire                weightFifo_6_pop_valid;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_6_pop_payload_1_2_2_15;
  wire                weightFifo_7_push_ready;
  wire                weightFifo_7_pop_valid;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_0_2_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_1_2_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_0_2_2_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_0_2_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_1_2_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_0_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_1_15;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_0;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_1;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_2;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_3;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_4;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_5;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_6;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_7;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_8;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_9;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_10;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_11;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_12;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_13;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_14;
  wire       [7:0]    weightFifo_7_pop_payload_1_2_2_15;
  wire                window_videoIn_ready;
  wire                window_videoOut_valid;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_payload_frame_line_endOfLine;
  wire                window_videoOut_payload_frame_endOfFrame;
  wire                window_videoOut_payload_endOfPack;
  wire                window_videoOut_fork_io_input_ready;
  wire                window_videoOut_fork_io_outputs_0_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_0_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_0_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_0_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_1_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_1_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_1_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_1_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_2_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_2_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_2_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_2_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_3_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_3_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_3_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_3_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_4_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_4_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_4_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_4_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_5_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_5_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_5_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_5_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_6_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_6_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_6_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_6_payload_endOfPack;
  wire                window_videoOut_fork_io_outputs_7_valid;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_15;
  wire                window_videoOut_fork_io_outputs_7_payload_frame_line_endOfLine;
  wire                window_videoOut_fork_io_outputs_7_payload_frame_endOfFrame;
  wire                window_videoOut_fork_io_outputs_7_payload_endOfPack;
  wire                unit_0_inputs_ready;
  wire                unit_0_weights_ready;
  wire                unit_0_outputs_valid;
  wire       [23:0]   unit_0_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_0_outputs_payload_frame_line_pixel_1;
  wire                unit_0_outputs_payload_frame_line_endOfLine;
  wire                unit_0_outputs_payload_frame_endOfFrame;
  wire                unit_0_outputs_payload_endOfPack;
  wire                unit_1_inputs_ready;
  wire                unit_1_weights_ready;
  wire                unit_1_outputs_valid;
  wire       [23:0]   unit_1_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_1_outputs_payload_frame_line_pixel_1;
  wire                unit_1_outputs_payload_frame_line_endOfLine;
  wire                unit_1_outputs_payload_frame_endOfFrame;
  wire                unit_1_outputs_payload_endOfPack;
  wire                unit_2_inputs_ready;
  wire                unit_2_weights_ready;
  wire                unit_2_outputs_valid;
  wire       [23:0]   unit_2_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_2_outputs_payload_frame_line_pixel_1;
  wire                unit_2_outputs_payload_frame_line_endOfLine;
  wire                unit_2_outputs_payload_frame_endOfFrame;
  wire                unit_2_outputs_payload_endOfPack;
  wire                unit_3_inputs_ready;
  wire                unit_3_weights_ready;
  wire                unit_3_outputs_valid;
  wire       [23:0]   unit_3_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_3_outputs_payload_frame_line_pixel_1;
  wire                unit_3_outputs_payload_frame_line_endOfLine;
  wire                unit_3_outputs_payload_frame_endOfFrame;
  wire                unit_3_outputs_payload_endOfPack;
  wire                unit_4_inputs_ready;
  wire                unit_4_weights_ready;
  wire                unit_4_outputs_valid;
  wire       [23:0]   unit_4_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_4_outputs_payload_frame_line_pixel_1;
  wire                unit_4_outputs_payload_frame_line_endOfLine;
  wire                unit_4_outputs_payload_frame_endOfFrame;
  wire                unit_4_outputs_payload_endOfPack;
  wire                unit_5_inputs_ready;
  wire                unit_5_weights_ready;
  wire                unit_5_outputs_valid;
  wire       [23:0]   unit_5_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_5_outputs_payload_frame_line_pixel_1;
  wire                unit_5_outputs_payload_frame_line_endOfLine;
  wire                unit_5_outputs_payload_frame_endOfFrame;
  wire                unit_5_outputs_payload_endOfPack;
  wire                unit_6_inputs_ready;
  wire                unit_6_weights_ready;
  wire                unit_6_outputs_valid;
  wire       [23:0]   unit_6_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_6_outputs_payload_frame_line_pixel_1;
  wire                unit_6_outputs_payload_frame_line_endOfLine;
  wire                unit_6_outputs_payload_frame_endOfFrame;
  wire                unit_6_outputs_payload_endOfPack;
  wire                unit_7_inputs_ready;
  wire                unit_7_weights_ready;
  wire                unit_7_outputs_valid;
  wire       [23:0]   unit_7_outputs_payload_frame_line_pixel_0;
  wire       [23:0]   unit_7_outputs_payload_frame_line_pixel_1;
  wire                unit_7_outputs_payload_frame_line_endOfLine;
  wire                unit_7_outputs_payload_frame_endOfFrame;
  wire                unit_7_outputs_payload_endOfPack;
  wire                pool_videoIn_ready;
  wire                pool_videoOut_valid;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_0;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_1;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_2;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_3;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_4;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_5;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_6;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_7;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_8;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_9;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_10;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_11;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_12;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_13;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_14;
  wire       [7:0]    pool_videoOut_payload_frame_line_pixel_15;
  wire                pool_videoOut_payload_frame_line_endOfLine;
  wire                pool_videoOut_payload_frame_endOfFrame;
  wire                pool_videoOut_payload_endOfPack;
  wire                table_1_newTable_ready;
  wire                table_1_index_ready;
  wire                table_1_value_valid;
  wire       [7:0]    table_1_value_payload_0;
  wire       [7:0]    table_1_value_payload_1;
  wire       [7:0]    table_1_value_payload_2;
  wire       [7:0]    table_1_value_payload_3;
  wire       [7:0]    table_1_value_payload_4;
  wire       [7:0]    table_1_value_payload_5;
  wire       [7:0]    table_1_value_payload_6;
  wire       [7:0]    table_1_value_payload_7;
  wire       [7:0]    table_1_value_payload_8;
  wire       [7:0]    table_1_value_payload_9;
  wire       [7:0]    table_1_value_payload_10;
  wire       [7:0]    table_1_value_payload_11;
  wire       [7:0]    table_1_value_payload_12;
  wire       [7:0]    table_1_value_payload_13;
  wire       [7:0]    table_1_value_payload_14;
  wire       [7:0]    table_1_value_payload_15;
  wire                streamDemux_2_io_input_ready;
  wire                streamDemux_2_io_outputs_0_valid;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_1_valid;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_2_valid;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_2_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_3_valid;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_3_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_4_valid;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_4_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_5_valid;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_5_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_6_valid;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_6_payload_1_2_2_15;
  wire                streamDemux_2_io_outputs_7_valid;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_0_2_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_0_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_1_2_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_0_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_1_15;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_0;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_1;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_2;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_3;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_4;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_5;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_6;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_7;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_8;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_9;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_10;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_11;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_12;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_13;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_14;
  wire       [7:0]    streamDemux_2_io_outputs_7_payload_1_2_2_15;
  wire                eventM2sPipes_9_eventIn_ready;
  wire                eventM2sPipes_9_eventOut_valid;
  wire                eventM2sPipes_9_CEs_0;
  wire                eventM2sPipes_9_CEs_1;
  wire                eventM2sPipes_9_CEs_2;
  wire                eventM2sPipes_9_CEs_3;
  wire                eventM2sPipes_9_CEs_4;
  wire                eventM2sPipes_9_CEs_5;
  wire       [7:0]    scalerINT16_16_dout;
  wire       [7:0]    scalerINT16_17_dout;
  wire       [7:0]    scalerINT16_18_dout;
  wire       [7:0]    scalerINT16_19_dout;
  wire       [7:0]    scalerINT16_20_dout;
  wire       [7:0]    scalerINT16_21_dout;
  wire       [7:0]    scalerINT16_22_dout;
  wire       [7:0]    scalerINT16_23_dout;
  wire       [7:0]    scalerINT16_24_dout;
  wire       [7:0]    scalerINT16_25_dout;
  wire       [7:0]    scalerINT16_26_dout;
  wire       [7:0]    scalerINT16_27_dout;
  wire       [7:0]    scalerINT16_28_dout;
  wire       [7:0]    scalerINT16_29_dout;
  wire       [7:0]    scalerINT16_30_dout;
  wire       [7:0]    scalerINT16_31_dout;
  wire                streamDemux_3_io_input_ready;
  wire                streamDemux_3_io_outputs_0_valid;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_0;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_1;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_2;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_3;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_4;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_5;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_6;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_7;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_8;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_9;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_10;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_11;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_12;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_13;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_14;
  wire       [7:0]    streamDemux_3_io_outputs_0_payload_frame_line_pixel_15;
  wire                streamDemux_3_io_outputs_0_payload_frame_line_endOfLine;
  wire                streamDemux_3_io_outputs_0_payload_frame_endOfFrame;
  wire                streamDemux_3_io_outputs_0_payload_endOfPack;
  wire                streamDemux_3_io_outputs_1_valid;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_0;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_1;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_2;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_3;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_4;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_5;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_6;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_7;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_8;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_9;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_10;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_11;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_12;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_13;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_14;
  wire       [7:0]    streamDemux_3_io_outputs_1_payload_frame_line_pixel_15;
  wire                streamDemux_3_io_outputs_1_payload_frame_line_endOfLine;
  wire                streamDemux_3_io_outputs_1_payload_frame_endOfFrame;
  wire                streamDemux_3_io_outputs_1_payload_endOfPack;
  wire                streamMux_1_io_inputs_0_ready;
  wire                streamMux_1_io_inputs_1_ready;
  wire                streamMux_1_io_output_valid;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_0;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_1;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_2;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_3;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_4;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_5;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_6;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_7;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_8;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_9;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_10;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_11;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_12;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_13;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_14;
  wire       [7:0]    streamMux_1_io_output_payload_frame_line_pixel_15;
  wire                streamMux_1_io_output_payload_frame_line_endOfLine;
  wire                streamMux_1_io_output_payload_frame_endOfFrame;
  wire                streamMux_1_io_output_payload_endOfPack;
  wire       [8:0]    tmp_tmp_when_Utils_l503_3;
  wire       [0:0]    tmp_tmp_when_Utils_l503_3_1;
  wire       [8:0]    tmp_tmp_when_Utils_l503_6;
  wire       [0:0]    tmp_tmp_when_Utils_l503_6_1;
  wire       [7:0]    tmp_tmp_inputVideo_payload_endOfPack_1;
  wire       [0:0]    tmp_tmp_inputVideo_payload_endOfPack_1_1;
  wire       [2:0]    tmp_tmp_io_select_1;
  wire       [0:0]    tmp_tmp_io_select_1_1;
  wire       [4:0]    tmp_tmp_weights_ready_1;
  wire       [0:0]    tmp_tmp_weights_ready_1_1;
  wire       [2047:0] tmp_tmp_weightsAdapted_payload_0_0_0_0;
  wire       [3:0]    tmp_tmp_funcTable_ready_1;
  wire       [0:0]    tmp_tmp_funcTable_ready_1_1;
  reg        [7:0]    tmp_tableAdapted_payload_1;
  wire                inputChannelSpilt_valid;
  wire                inputChannelSpilt_ready;
  wire       [7:0]    inputChannelSpilt_payload_0;
  wire       [7:0]    inputChannelSpilt_payload_1;
  wire       [7:0]    inputChannelSpilt_payload_2;
  wire       [7:0]    inputChannelSpilt_payload_3;
  wire       [7:0]    inputChannelSpilt_payload_4;
  wire       [7:0]    inputChannelSpilt_payload_5;
  wire       [7:0]    inputChannelSpilt_payload_6;
  wire       [7:0]    inputChannelSpilt_payload_7;
  wire       [7:0]    inputChannelSpilt_payload_8;
  wire       [7:0]    inputChannelSpilt_payload_9;
  wire       [7:0]    inputChannelSpilt_payload_10;
  wire       [7:0]    inputChannelSpilt_payload_11;
  wire       [7:0]    inputChannelSpilt_payload_12;
  wire       [7:0]    inputChannelSpilt_payload_13;
  wire       [7:0]    inputChannelSpilt_payload_14;
  wire       [7:0]    inputChannelSpilt_payload_15;
  wire       [127:0]  tmp_inputChannelSpilt_payload_0;
  wire                inputChannelSpilt_translated_valid;
  reg                 inputChannelSpilt_translated_ready;
  wire       [7:0]    inputChannelSpilt_translated_payload_0;
  wire       [7:0]    inputChannelSpilt_translated_payload_1;
  wire       [7:0]    inputChannelSpilt_translated_payload_2;
  wire       [7:0]    inputChannelSpilt_translated_payload_3;
  wire       [7:0]    inputChannelSpilt_translated_payload_4;
  wire       [7:0]    inputChannelSpilt_translated_payload_5;
  wire       [7:0]    inputChannelSpilt_translated_payload_6;
  wire       [7:0]    inputChannelSpilt_translated_payload_7;
  wire       [7:0]    inputChannelSpilt_translated_payload_8;
  wire       [7:0]    inputChannelSpilt_translated_payload_9;
  wire       [7:0]    inputChannelSpilt_translated_payload_10;
  wire       [7:0]    inputChannelSpilt_translated_payload_11;
  wire       [7:0]    inputChannelSpilt_translated_payload_12;
  wire       [7:0]    inputChannelSpilt_translated_payload_13;
  wire       [7:0]    inputChannelSpilt_translated_payload_14;
  wire       [7:0]    inputChannelSpilt_translated_payload_15;
  wire                inputChannelSpilt_translated_m2sPipe_valid;
  wire                inputChannelSpilt_translated_m2sPipe_ready;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_0;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_1;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_2;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_3;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_4;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_5;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_6;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_7;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_8;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_9;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_10;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_11;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_12;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_13;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_14;
  wire       [7:0]    inputChannelSpilt_translated_m2sPipe_payload_15;
  reg                 inputChannelSpilt_translated_rValid;
  reg        [7:0]    inputChannelSpilt_translated_rData_0;
  reg        [7:0]    inputChannelSpilt_translated_rData_1;
  reg        [7:0]    inputChannelSpilt_translated_rData_2;
  reg        [7:0]    inputChannelSpilt_translated_rData_3;
  reg        [7:0]    inputChannelSpilt_translated_rData_4;
  reg        [7:0]    inputChannelSpilt_translated_rData_5;
  reg        [7:0]    inputChannelSpilt_translated_rData_6;
  reg        [7:0]    inputChannelSpilt_translated_rData_7;
  reg        [7:0]    inputChannelSpilt_translated_rData_8;
  reg        [7:0]    inputChannelSpilt_translated_rData_9;
  reg        [7:0]    inputChannelSpilt_translated_rData_10;
  reg        [7:0]    inputChannelSpilt_translated_rData_11;
  reg        [7:0]    inputChannelSpilt_translated_rData_12;
  reg        [7:0]    inputChannelSpilt_translated_rData_13;
  reg        [7:0]    inputChannelSpilt_translated_rData_14;
  reg        [7:0]    inputChannelSpilt_translated_rData_15;
  wire                when_Stream_l342;
  wire                inputChannelSpilt_translated_m2sPipe_fire;
  wire                tmp_when_Utils_l503;
  wire                tmp_when_Utils_l503_1;
  reg                 tmp_when_Utils_l503_2;
  reg        [8:0]    tmp_when_Utils_l503_3;
  reg        [8:0]    tmp_when_Utils_l503_4;
  wire                when_Utils_l503;
  reg                 tmp_when_Utils_l503_5;
  reg        [8:0]    tmp_when_Utils_l503_6;
  reg        [8:0]    tmp_when_Utils_l503_7;
  wire                when_Utils_l503_1;
  reg                 tmp_inputVideo_payload_endOfPack;
  reg        [7:0]    tmp_inputVideo_payload_endOfPack_1;
  reg        [7:0]    tmp_inputVideo_payload_endOfPack_2;
  wire                inputVideo_valid;
  wire                inputVideo_ready;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_0;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_1;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_2;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_3;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_4;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_5;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_6;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_7;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_8;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_9;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_10;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_11;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_12;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_13;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_14;
  wire       [7:0]    inputVideo_payload_frame_line_pixel_15;
  wire                inputVideo_payload_frame_line_endOfLine;
  wire                inputVideo_payload_frame_endOfFrame;
  wire                inputVideo_payload_endOfPack;
  wire                weightsAdapted_valid;
  wire                weightsAdapted_ready;
  wire       [7:0]    weightsAdapted_payload_0_0_0_0;
  wire       [7:0]    weightsAdapted_payload_0_0_0_1;
  wire       [7:0]    weightsAdapted_payload_0_0_0_2;
  wire       [7:0]    weightsAdapted_payload_0_0_0_3;
  wire       [7:0]    weightsAdapted_payload_0_0_0_4;
  wire       [7:0]    weightsAdapted_payload_0_0_0_5;
  wire       [7:0]    weightsAdapted_payload_0_0_0_6;
  wire       [7:0]    weightsAdapted_payload_0_0_0_7;
  wire       [7:0]    weightsAdapted_payload_0_0_0_8;
  wire       [7:0]    weightsAdapted_payload_0_0_0_9;
  wire       [7:0]    weightsAdapted_payload_0_0_0_10;
  wire       [7:0]    weightsAdapted_payload_0_0_0_11;
  wire       [7:0]    weightsAdapted_payload_0_0_0_12;
  wire       [7:0]    weightsAdapted_payload_0_0_0_13;
  wire       [7:0]    weightsAdapted_payload_0_0_0_14;
  wire       [7:0]    weightsAdapted_payload_0_0_0_15;
  wire       [7:0]    weightsAdapted_payload_0_0_1_0;
  wire       [7:0]    weightsAdapted_payload_0_0_1_1;
  wire       [7:0]    weightsAdapted_payload_0_0_1_2;
  wire       [7:0]    weightsAdapted_payload_0_0_1_3;
  wire       [7:0]    weightsAdapted_payload_0_0_1_4;
  wire       [7:0]    weightsAdapted_payload_0_0_1_5;
  wire       [7:0]    weightsAdapted_payload_0_0_1_6;
  wire       [7:0]    weightsAdapted_payload_0_0_1_7;
  wire       [7:0]    weightsAdapted_payload_0_0_1_8;
  wire       [7:0]    weightsAdapted_payload_0_0_1_9;
  wire       [7:0]    weightsAdapted_payload_0_0_1_10;
  wire       [7:0]    weightsAdapted_payload_0_0_1_11;
  wire       [7:0]    weightsAdapted_payload_0_0_1_12;
  wire       [7:0]    weightsAdapted_payload_0_0_1_13;
  wire       [7:0]    weightsAdapted_payload_0_0_1_14;
  wire       [7:0]    weightsAdapted_payload_0_0_1_15;
  wire       [7:0]    weightsAdapted_payload_0_0_2_0;
  wire       [7:0]    weightsAdapted_payload_0_0_2_1;
  wire       [7:0]    weightsAdapted_payload_0_0_2_2;
  wire       [7:0]    weightsAdapted_payload_0_0_2_3;
  wire       [7:0]    weightsAdapted_payload_0_0_2_4;
  wire       [7:0]    weightsAdapted_payload_0_0_2_5;
  wire       [7:0]    weightsAdapted_payload_0_0_2_6;
  wire       [7:0]    weightsAdapted_payload_0_0_2_7;
  wire       [7:0]    weightsAdapted_payload_0_0_2_8;
  wire       [7:0]    weightsAdapted_payload_0_0_2_9;
  wire       [7:0]    weightsAdapted_payload_0_0_2_10;
  wire       [7:0]    weightsAdapted_payload_0_0_2_11;
  wire       [7:0]    weightsAdapted_payload_0_0_2_12;
  wire       [7:0]    weightsAdapted_payload_0_0_2_13;
  wire       [7:0]    weightsAdapted_payload_0_0_2_14;
  wire       [7:0]    weightsAdapted_payload_0_0_2_15;
  wire       [7:0]    weightsAdapted_payload_0_1_0_0;
  wire       [7:0]    weightsAdapted_payload_0_1_0_1;
  wire       [7:0]    weightsAdapted_payload_0_1_0_2;
  wire       [7:0]    weightsAdapted_payload_0_1_0_3;
  wire       [7:0]    weightsAdapted_payload_0_1_0_4;
  wire       [7:0]    weightsAdapted_payload_0_1_0_5;
  wire       [7:0]    weightsAdapted_payload_0_1_0_6;
  wire       [7:0]    weightsAdapted_payload_0_1_0_7;
  wire       [7:0]    weightsAdapted_payload_0_1_0_8;
  wire       [7:0]    weightsAdapted_payload_0_1_0_9;
  wire       [7:0]    weightsAdapted_payload_0_1_0_10;
  wire       [7:0]    weightsAdapted_payload_0_1_0_11;
  wire       [7:0]    weightsAdapted_payload_0_1_0_12;
  wire       [7:0]    weightsAdapted_payload_0_1_0_13;
  wire       [7:0]    weightsAdapted_payload_0_1_0_14;
  wire       [7:0]    weightsAdapted_payload_0_1_0_15;
  wire       [7:0]    weightsAdapted_payload_0_1_1_0;
  wire       [7:0]    weightsAdapted_payload_0_1_1_1;
  wire       [7:0]    weightsAdapted_payload_0_1_1_2;
  wire       [7:0]    weightsAdapted_payload_0_1_1_3;
  wire       [7:0]    weightsAdapted_payload_0_1_1_4;
  wire       [7:0]    weightsAdapted_payload_0_1_1_5;
  wire       [7:0]    weightsAdapted_payload_0_1_1_6;
  wire       [7:0]    weightsAdapted_payload_0_1_1_7;
  wire       [7:0]    weightsAdapted_payload_0_1_1_8;
  wire       [7:0]    weightsAdapted_payload_0_1_1_9;
  wire       [7:0]    weightsAdapted_payload_0_1_1_10;
  wire       [7:0]    weightsAdapted_payload_0_1_1_11;
  wire       [7:0]    weightsAdapted_payload_0_1_1_12;
  wire       [7:0]    weightsAdapted_payload_0_1_1_13;
  wire       [7:0]    weightsAdapted_payload_0_1_1_14;
  wire       [7:0]    weightsAdapted_payload_0_1_1_15;
  wire       [7:0]    weightsAdapted_payload_0_1_2_0;
  wire       [7:0]    weightsAdapted_payload_0_1_2_1;
  wire       [7:0]    weightsAdapted_payload_0_1_2_2;
  wire       [7:0]    weightsAdapted_payload_0_1_2_3;
  wire       [7:0]    weightsAdapted_payload_0_1_2_4;
  wire       [7:0]    weightsAdapted_payload_0_1_2_5;
  wire       [7:0]    weightsAdapted_payload_0_1_2_6;
  wire       [7:0]    weightsAdapted_payload_0_1_2_7;
  wire       [7:0]    weightsAdapted_payload_0_1_2_8;
  wire       [7:0]    weightsAdapted_payload_0_1_2_9;
  wire       [7:0]    weightsAdapted_payload_0_1_2_10;
  wire       [7:0]    weightsAdapted_payload_0_1_2_11;
  wire       [7:0]    weightsAdapted_payload_0_1_2_12;
  wire       [7:0]    weightsAdapted_payload_0_1_2_13;
  wire       [7:0]    weightsAdapted_payload_0_1_2_14;
  wire       [7:0]    weightsAdapted_payload_0_1_2_15;
  wire       [7:0]    weightsAdapted_payload_0_2_0_0;
  wire       [7:0]    weightsAdapted_payload_0_2_0_1;
  wire       [7:0]    weightsAdapted_payload_0_2_0_2;
  wire       [7:0]    weightsAdapted_payload_0_2_0_3;
  wire       [7:0]    weightsAdapted_payload_0_2_0_4;
  wire       [7:0]    weightsAdapted_payload_0_2_0_5;
  wire       [7:0]    weightsAdapted_payload_0_2_0_6;
  wire       [7:0]    weightsAdapted_payload_0_2_0_7;
  wire       [7:0]    weightsAdapted_payload_0_2_0_8;
  wire       [7:0]    weightsAdapted_payload_0_2_0_9;
  wire       [7:0]    weightsAdapted_payload_0_2_0_10;
  wire       [7:0]    weightsAdapted_payload_0_2_0_11;
  wire       [7:0]    weightsAdapted_payload_0_2_0_12;
  wire       [7:0]    weightsAdapted_payload_0_2_0_13;
  wire       [7:0]    weightsAdapted_payload_0_2_0_14;
  wire       [7:0]    weightsAdapted_payload_0_2_0_15;
  wire       [7:0]    weightsAdapted_payload_0_2_1_0;
  wire       [7:0]    weightsAdapted_payload_0_2_1_1;
  wire       [7:0]    weightsAdapted_payload_0_2_1_2;
  wire       [7:0]    weightsAdapted_payload_0_2_1_3;
  wire       [7:0]    weightsAdapted_payload_0_2_1_4;
  wire       [7:0]    weightsAdapted_payload_0_2_1_5;
  wire       [7:0]    weightsAdapted_payload_0_2_1_6;
  wire       [7:0]    weightsAdapted_payload_0_2_1_7;
  wire       [7:0]    weightsAdapted_payload_0_2_1_8;
  wire       [7:0]    weightsAdapted_payload_0_2_1_9;
  wire       [7:0]    weightsAdapted_payload_0_2_1_10;
  wire       [7:0]    weightsAdapted_payload_0_2_1_11;
  wire       [7:0]    weightsAdapted_payload_0_2_1_12;
  wire       [7:0]    weightsAdapted_payload_0_2_1_13;
  wire       [7:0]    weightsAdapted_payload_0_2_1_14;
  wire       [7:0]    weightsAdapted_payload_0_2_1_15;
  wire       [7:0]    weightsAdapted_payload_0_2_2_0;
  wire       [7:0]    weightsAdapted_payload_0_2_2_1;
  wire       [7:0]    weightsAdapted_payload_0_2_2_2;
  wire       [7:0]    weightsAdapted_payload_0_2_2_3;
  wire       [7:0]    weightsAdapted_payload_0_2_2_4;
  wire       [7:0]    weightsAdapted_payload_0_2_2_5;
  wire       [7:0]    weightsAdapted_payload_0_2_2_6;
  wire       [7:0]    weightsAdapted_payload_0_2_2_7;
  wire       [7:0]    weightsAdapted_payload_0_2_2_8;
  wire       [7:0]    weightsAdapted_payload_0_2_2_9;
  wire       [7:0]    weightsAdapted_payload_0_2_2_10;
  wire       [7:0]    weightsAdapted_payload_0_2_2_11;
  wire       [7:0]    weightsAdapted_payload_0_2_2_12;
  wire       [7:0]    weightsAdapted_payload_0_2_2_13;
  wire       [7:0]    weightsAdapted_payload_0_2_2_14;
  wire       [7:0]    weightsAdapted_payload_0_2_2_15;
  wire       [7:0]    weightsAdapted_payload_1_0_0_0;
  wire       [7:0]    weightsAdapted_payload_1_0_0_1;
  wire       [7:0]    weightsAdapted_payload_1_0_0_2;
  wire       [7:0]    weightsAdapted_payload_1_0_0_3;
  wire       [7:0]    weightsAdapted_payload_1_0_0_4;
  wire       [7:0]    weightsAdapted_payload_1_0_0_5;
  wire       [7:0]    weightsAdapted_payload_1_0_0_6;
  wire       [7:0]    weightsAdapted_payload_1_0_0_7;
  wire       [7:0]    weightsAdapted_payload_1_0_0_8;
  wire       [7:0]    weightsAdapted_payload_1_0_0_9;
  wire       [7:0]    weightsAdapted_payload_1_0_0_10;
  wire       [7:0]    weightsAdapted_payload_1_0_0_11;
  wire       [7:0]    weightsAdapted_payload_1_0_0_12;
  wire       [7:0]    weightsAdapted_payload_1_0_0_13;
  wire       [7:0]    weightsAdapted_payload_1_0_0_14;
  wire       [7:0]    weightsAdapted_payload_1_0_0_15;
  wire       [7:0]    weightsAdapted_payload_1_0_1_0;
  wire       [7:0]    weightsAdapted_payload_1_0_1_1;
  wire       [7:0]    weightsAdapted_payload_1_0_1_2;
  wire       [7:0]    weightsAdapted_payload_1_0_1_3;
  wire       [7:0]    weightsAdapted_payload_1_0_1_4;
  wire       [7:0]    weightsAdapted_payload_1_0_1_5;
  wire       [7:0]    weightsAdapted_payload_1_0_1_6;
  wire       [7:0]    weightsAdapted_payload_1_0_1_7;
  wire       [7:0]    weightsAdapted_payload_1_0_1_8;
  wire       [7:0]    weightsAdapted_payload_1_0_1_9;
  wire       [7:0]    weightsAdapted_payload_1_0_1_10;
  wire       [7:0]    weightsAdapted_payload_1_0_1_11;
  wire       [7:0]    weightsAdapted_payload_1_0_1_12;
  wire       [7:0]    weightsAdapted_payload_1_0_1_13;
  wire       [7:0]    weightsAdapted_payload_1_0_1_14;
  wire       [7:0]    weightsAdapted_payload_1_0_1_15;
  wire       [7:0]    weightsAdapted_payload_1_0_2_0;
  wire       [7:0]    weightsAdapted_payload_1_0_2_1;
  wire       [7:0]    weightsAdapted_payload_1_0_2_2;
  wire       [7:0]    weightsAdapted_payload_1_0_2_3;
  wire       [7:0]    weightsAdapted_payload_1_0_2_4;
  wire       [7:0]    weightsAdapted_payload_1_0_2_5;
  wire       [7:0]    weightsAdapted_payload_1_0_2_6;
  wire       [7:0]    weightsAdapted_payload_1_0_2_7;
  wire       [7:0]    weightsAdapted_payload_1_0_2_8;
  wire       [7:0]    weightsAdapted_payload_1_0_2_9;
  wire       [7:0]    weightsAdapted_payload_1_0_2_10;
  wire       [7:0]    weightsAdapted_payload_1_0_2_11;
  wire       [7:0]    weightsAdapted_payload_1_0_2_12;
  wire       [7:0]    weightsAdapted_payload_1_0_2_13;
  wire       [7:0]    weightsAdapted_payload_1_0_2_14;
  wire       [7:0]    weightsAdapted_payload_1_0_2_15;
  wire       [7:0]    weightsAdapted_payload_1_1_0_0;
  wire       [7:0]    weightsAdapted_payload_1_1_0_1;
  wire       [7:0]    weightsAdapted_payload_1_1_0_2;
  wire       [7:0]    weightsAdapted_payload_1_1_0_3;
  wire       [7:0]    weightsAdapted_payload_1_1_0_4;
  wire       [7:0]    weightsAdapted_payload_1_1_0_5;
  wire       [7:0]    weightsAdapted_payload_1_1_0_6;
  wire       [7:0]    weightsAdapted_payload_1_1_0_7;
  wire       [7:0]    weightsAdapted_payload_1_1_0_8;
  wire       [7:0]    weightsAdapted_payload_1_1_0_9;
  wire       [7:0]    weightsAdapted_payload_1_1_0_10;
  wire       [7:0]    weightsAdapted_payload_1_1_0_11;
  wire       [7:0]    weightsAdapted_payload_1_1_0_12;
  wire       [7:0]    weightsAdapted_payload_1_1_0_13;
  wire       [7:0]    weightsAdapted_payload_1_1_0_14;
  wire       [7:0]    weightsAdapted_payload_1_1_0_15;
  wire       [7:0]    weightsAdapted_payload_1_1_1_0;
  wire       [7:0]    weightsAdapted_payload_1_1_1_1;
  wire       [7:0]    weightsAdapted_payload_1_1_1_2;
  wire       [7:0]    weightsAdapted_payload_1_1_1_3;
  wire       [7:0]    weightsAdapted_payload_1_1_1_4;
  wire       [7:0]    weightsAdapted_payload_1_1_1_5;
  wire       [7:0]    weightsAdapted_payload_1_1_1_6;
  wire       [7:0]    weightsAdapted_payload_1_1_1_7;
  wire       [7:0]    weightsAdapted_payload_1_1_1_8;
  wire       [7:0]    weightsAdapted_payload_1_1_1_9;
  wire       [7:0]    weightsAdapted_payload_1_1_1_10;
  wire       [7:0]    weightsAdapted_payload_1_1_1_11;
  wire       [7:0]    weightsAdapted_payload_1_1_1_12;
  wire       [7:0]    weightsAdapted_payload_1_1_1_13;
  wire       [7:0]    weightsAdapted_payload_1_1_1_14;
  wire       [7:0]    weightsAdapted_payload_1_1_1_15;
  wire       [7:0]    weightsAdapted_payload_1_1_2_0;
  wire       [7:0]    weightsAdapted_payload_1_1_2_1;
  wire       [7:0]    weightsAdapted_payload_1_1_2_2;
  wire       [7:0]    weightsAdapted_payload_1_1_2_3;
  wire       [7:0]    weightsAdapted_payload_1_1_2_4;
  wire       [7:0]    weightsAdapted_payload_1_1_2_5;
  wire       [7:0]    weightsAdapted_payload_1_1_2_6;
  wire       [7:0]    weightsAdapted_payload_1_1_2_7;
  wire       [7:0]    weightsAdapted_payload_1_1_2_8;
  wire       [7:0]    weightsAdapted_payload_1_1_2_9;
  wire       [7:0]    weightsAdapted_payload_1_1_2_10;
  wire       [7:0]    weightsAdapted_payload_1_1_2_11;
  wire       [7:0]    weightsAdapted_payload_1_1_2_12;
  wire       [7:0]    weightsAdapted_payload_1_1_2_13;
  wire       [7:0]    weightsAdapted_payload_1_1_2_14;
  wire       [7:0]    weightsAdapted_payload_1_1_2_15;
  wire       [7:0]    weightsAdapted_payload_1_2_0_0;
  wire       [7:0]    weightsAdapted_payload_1_2_0_1;
  wire       [7:0]    weightsAdapted_payload_1_2_0_2;
  wire       [7:0]    weightsAdapted_payload_1_2_0_3;
  wire       [7:0]    weightsAdapted_payload_1_2_0_4;
  wire       [7:0]    weightsAdapted_payload_1_2_0_5;
  wire       [7:0]    weightsAdapted_payload_1_2_0_6;
  wire       [7:0]    weightsAdapted_payload_1_2_0_7;
  wire       [7:0]    weightsAdapted_payload_1_2_0_8;
  wire       [7:0]    weightsAdapted_payload_1_2_0_9;
  wire       [7:0]    weightsAdapted_payload_1_2_0_10;
  wire       [7:0]    weightsAdapted_payload_1_2_0_11;
  wire       [7:0]    weightsAdapted_payload_1_2_0_12;
  wire       [7:0]    weightsAdapted_payload_1_2_0_13;
  wire       [7:0]    weightsAdapted_payload_1_2_0_14;
  wire       [7:0]    weightsAdapted_payload_1_2_0_15;
  wire       [7:0]    weightsAdapted_payload_1_2_1_0;
  wire       [7:0]    weightsAdapted_payload_1_2_1_1;
  wire       [7:0]    weightsAdapted_payload_1_2_1_2;
  wire       [7:0]    weightsAdapted_payload_1_2_1_3;
  wire       [7:0]    weightsAdapted_payload_1_2_1_4;
  wire       [7:0]    weightsAdapted_payload_1_2_1_5;
  wire       [7:0]    weightsAdapted_payload_1_2_1_6;
  wire       [7:0]    weightsAdapted_payload_1_2_1_7;
  wire       [7:0]    weightsAdapted_payload_1_2_1_8;
  wire       [7:0]    weightsAdapted_payload_1_2_1_9;
  wire       [7:0]    weightsAdapted_payload_1_2_1_10;
  wire       [7:0]    weightsAdapted_payload_1_2_1_11;
  wire       [7:0]    weightsAdapted_payload_1_2_1_12;
  wire       [7:0]    weightsAdapted_payload_1_2_1_13;
  wire       [7:0]    weightsAdapted_payload_1_2_1_14;
  wire       [7:0]    weightsAdapted_payload_1_2_1_15;
  wire       [7:0]    weightsAdapted_payload_1_2_2_0;
  wire       [7:0]    weightsAdapted_payload_1_2_2_1;
  wire       [7:0]    weightsAdapted_payload_1_2_2_2;
  wire       [7:0]    weightsAdapted_payload_1_2_2_3;
  wire       [7:0]    weightsAdapted_payload_1_2_2_4;
  wire       [7:0]    weightsAdapted_payload_1_2_2_5;
  wire       [7:0]    weightsAdapted_payload_1_2_2_6;
  wire       [7:0]    weightsAdapted_payload_1_2_2_7;
  wire       [7:0]    weightsAdapted_payload_1_2_2_8;
  wire       [7:0]    weightsAdapted_payload_1_2_2_9;
  wire       [7:0]    weightsAdapted_payload_1_2_2_10;
  wire       [7:0]    weightsAdapted_payload_1_2_2_11;
  wire       [7:0]    weightsAdapted_payload_1_2_2_12;
  wire       [7:0]    weightsAdapted_payload_1_2_2_13;
  wire       [7:0]    weightsAdapted_payload_1_2_2_14;
  wire       [7:0]    weightsAdapted_payload_1_2_2_15;
  reg                 tmp_io_select;
  reg        [2:0]    tmp_io_select_1;
  reg        [2:0]    tmp_io_select_2;
  wire                weightsAdapted_fire;
  wire                weights_fire;
  reg                 tmp_weights_ready;
  reg        [4:0]    tmp_weights_ready_1;
  reg        [4:0]    tmp_weights_ready_2;
  wire                tmp_weights_ready_3;
  wire                tmp_1;
  reg        [2175:0] tmp_weightsAdapted_payload_0_0_0_0;
  wire                weights_fire_1;
  wire       [2303:0] tmp_weightsAdapted_payload_0_0_0_0_1;
  wire       [1151:0] tmp_weightsAdapted_payload_0_0_0_0_2;
  wire       [383:0]  tmp_weightsAdapted_payload_0_0_0_0_3;
  wire       [127:0]  tmp_weightsAdapted_payload_0_0_0_0_4;
  wire       [127:0]  tmp_weightsAdapted_payload_0_0_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_0_0_2_0;
  wire       [383:0]  tmp_weightsAdapted_payload_0_1_0_0;
  wire       [127:0]  tmp_weightsAdapted_payload_0_1_0_0_1;
  wire       [127:0]  tmp_weightsAdapted_payload_0_1_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_0_1_2_0;
  wire       [383:0]  tmp_weightsAdapted_payload_0_2_0_0;
  wire       [127:0]  tmp_weightsAdapted_payload_0_2_0_0_1;
  wire       [127:0]  tmp_weightsAdapted_payload_0_2_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_0_2_2_0;
  wire       [1151:0] tmp_weightsAdapted_payload_1_0_0_0;
  wire       [383:0]  tmp_weightsAdapted_payload_1_0_0_0_1;
  wire       [127:0]  tmp_weightsAdapted_payload_1_0_0_0_2;
  wire       [127:0]  tmp_weightsAdapted_payload_1_0_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_1_0_2_0;
  wire       [383:0]  tmp_weightsAdapted_payload_1_1_0_0;
  wire       [127:0]  tmp_weightsAdapted_payload_1_1_0_0_1;
  wire       [127:0]  tmp_weightsAdapted_payload_1_1_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_1_1_2_0;
  wire       [383:0]  tmp_weightsAdapted_payload_1_2_0_0;
  wire       [127:0]  tmp_weightsAdapted_payload_1_2_0_0_1;
  wire       [127:0]  tmp_weightsAdapted_payload_1_2_1_0;
  wire       [127:0]  tmp_weightsAdapted_payload_1_2_2_0;
  wire                accOutputs_0_valid;
  wire                accOutputs_0_ready;
  wire       [23:0]   accOutputs_0_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_0_payload_frame_line_pixel_1;
  wire                accOutputs_0_payload_frame_line_endOfLine;
  wire                accOutputs_0_payload_frame_endOfFrame;
  wire                accOutputs_0_payload_endOfPack;
  wire                accOutputs_1_valid;
  wire                accOutputs_1_ready;
  wire       [23:0]   accOutputs_1_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_1_payload_frame_line_pixel_1;
  wire                accOutputs_1_payload_frame_line_endOfLine;
  wire                accOutputs_1_payload_frame_endOfFrame;
  wire                accOutputs_1_payload_endOfPack;
  wire                accOutputs_2_valid;
  wire                accOutputs_2_ready;
  wire       [23:0]   accOutputs_2_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_2_payload_frame_line_pixel_1;
  wire                accOutputs_2_payload_frame_line_endOfLine;
  wire                accOutputs_2_payload_frame_endOfFrame;
  wire                accOutputs_2_payload_endOfPack;
  wire                accOutputs_3_valid;
  wire                accOutputs_3_ready;
  wire       [23:0]   accOutputs_3_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_3_payload_frame_line_pixel_1;
  wire                accOutputs_3_payload_frame_line_endOfLine;
  wire                accOutputs_3_payload_frame_endOfFrame;
  wire                accOutputs_3_payload_endOfPack;
  wire                accOutputs_4_valid;
  wire                accOutputs_4_ready;
  wire       [23:0]   accOutputs_4_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_4_payload_frame_line_pixel_1;
  wire                accOutputs_4_payload_frame_line_endOfLine;
  wire                accOutputs_4_payload_frame_endOfFrame;
  wire                accOutputs_4_payload_endOfPack;
  wire                accOutputs_5_valid;
  wire                accOutputs_5_ready;
  wire       [23:0]   accOutputs_5_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_5_payload_frame_line_pixel_1;
  wire                accOutputs_5_payload_frame_line_endOfLine;
  wire                accOutputs_5_payload_frame_endOfFrame;
  wire                accOutputs_5_payload_endOfPack;
  wire                accOutputs_6_valid;
  wire                accOutputs_6_ready;
  wire       [23:0]   accOutputs_6_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_6_payload_frame_line_pixel_1;
  wire                accOutputs_6_payload_frame_line_endOfLine;
  wire                accOutputs_6_payload_frame_endOfFrame;
  wire                accOutputs_6_payload_endOfPack;
  wire                accOutputs_7_valid;
  wire                accOutputs_7_ready;
  wire       [23:0]   accOutputs_7_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputs_7_payload_frame_line_pixel_1;
  wire                accOutputs_7_payload_frame_line_endOfLine;
  wire                accOutputs_7_payload_frame_endOfFrame;
  wire                accOutputs_7_payload_endOfPack;
  wire                accOutputsJoin_valid;
  wire                accOutputsJoin_ready;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_0;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_1;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_2;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_3;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_4;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_5;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_6;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_7;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_8;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_9;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_10;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_11;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_12;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_13;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_14;
  wire       [23:0]   accOutputsJoin_payload_frame_line_pixel_15;
  wire                accOutputsJoin_payload_frame_line_endOfLine;
  wire                accOutputsJoin_payload_frame_endOfFrame;
  wire                accOutputsJoin_payload_endOfPack;
  wire                tmp_accOutputs_0_ready;
  wire                tmp_accOutputs_0_ready_1;
  wire       [383:0]  tmp_accOutputsJoin_payload_frame_line_pixel_0;
  wire                postProcessOutputs_valid;
  wire                postProcessOutputs_ready;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_0;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_1;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_2;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_3;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_4;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_5;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_6;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_7;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_8;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_9;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_10;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_11;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_12;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_13;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_14;
  wire       [7:0]    postProcessOutputs_payload_frame_line_pixel_15;
  wire                postProcessOutputs_payload_frame_line_endOfLine;
  wire                postProcessOutputs_payload_frame_endOfFrame;
  wire                postProcessOutputs_payload_endOfPack;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame;
  reg                 tmp_postProcessOutputs_payload_endOfPack;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine_1;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame_1;
  reg                 tmp_postProcessOutputs_payload_endOfPack_1;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine_2;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame_2;
  reg                 tmp_postProcessOutputs_payload_endOfPack_2;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine_3;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame_3;
  reg                 tmp_postProcessOutputs_payload_endOfPack_3;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine_4;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame_4;
  reg                 tmp_postProcessOutputs_payload_endOfPack_4;
  reg                 tmp_postProcessOutputs_payload_frame_line_endOfLine_5;
  reg                 tmp_postProcessOutputs_payload_frame_endOfFrame_5;
  reg                 tmp_postProcessOutputs_payload_endOfPack_5;
  wire                tableAdapted_valid;
  wire                tableAdapted_ready;
  wire       [7:0]    tableAdapted_payload;
  wire                streamMux_1_io_output_translated_valid;
  wire                streamMux_1_io_output_translated_ready;
  wire       [7:0]    streamMux_1_io_output_translated_payload_0;
  wire       [7:0]    streamMux_1_io_output_translated_payload_1;
  wire       [7:0]    streamMux_1_io_output_translated_payload_2;
  wire       [7:0]    streamMux_1_io_output_translated_payload_3;
  wire       [7:0]    streamMux_1_io_output_translated_payload_4;
  wire       [7:0]    streamMux_1_io_output_translated_payload_5;
  wire       [7:0]    streamMux_1_io_output_translated_payload_6;
  wire       [7:0]    streamMux_1_io_output_translated_payload_7;
  wire       [7:0]    streamMux_1_io_output_translated_payload_8;
  wire       [7:0]    streamMux_1_io_output_translated_payload_9;
  wire       [7:0]    streamMux_1_io_output_translated_payload_10;
  wire       [7:0]    streamMux_1_io_output_translated_payload_11;
  wire       [7:0]    streamMux_1_io_output_translated_payload_12;
  wire       [7:0]    streamMux_1_io_output_translated_payload_13;
  wire       [7:0]    streamMux_1_io_output_translated_payload_14;
  wire       [7:0]    streamMux_1_io_output_translated_payload_15;
  wire                signalTrim_valid;
  wire                signalTrim_ready;
  wire       [7:0]    signalTrim_payload_0;
  wire       [7:0]    signalTrim_payload_1;
  wire       [7:0]    signalTrim_payload_2;
  wire       [7:0]    signalTrim_payload_3;
  wire       [7:0]    signalTrim_payload_4;
  wire       [7:0]    signalTrim_payload_5;
  wire       [7:0]    signalTrim_payload_6;
  wire       [7:0]    signalTrim_payload_7;
  wire       [7:0]    signalTrim_payload_8;
  wire       [7:0]    signalTrim_payload_9;
  wire       [7:0]    signalTrim_payload_10;
  wire       [7:0]    signalTrim_payload_11;
  wire       [7:0]    signalTrim_payload_12;
  wire       [7:0]    signalTrim_payload_13;
  wire       [7:0]    signalTrim_payload_14;
  wire       [7:0]    signalTrim_payload_15;
  wire       [127:0]  tmp_signalTrim_payload_0;
  wire                tableAdapted_fire;
  reg                 tmp_funcTable_ready;
  reg        [3:0]    tmp_funcTable_ready_1;
  reg        [3:0]    tmp_funcTable_ready_2;
  wire                tmp_funcTable_ready_3;
  wire       [127:0]  tmp_tableAdapted_payload;
  wire                table_1_value_transmuted_valid;
  wire                table_1_value_transmuted_ready;
  wire       [127:0]  table_1_value_transmuted_payload;

  assign tmp_tmp_when_Utils_l503_3_1 = tmp_when_Utils_l503_2;
  assign tmp_tmp_when_Utils_l503_3 = {8'd0, tmp_tmp_when_Utils_l503_3_1};
  assign tmp_tmp_when_Utils_l503_6_1 = tmp_when_Utils_l503_5;
  assign tmp_tmp_when_Utils_l503_6 = {8'd0, tmp_tmp_when_Utils_l503_6_1};
  assign tmp_tmp_inputVideo_payload_endOfPack_1_1 = tmp_inputVideo_payload_endOfPack;
  assign tmp_tmp_inputVideo_payload_endOfPack_1 = {7'd0, tmp_tmp_inputVideo_payload_endOfPack_1_1};
  assign tmp_tmp_io_select_1_1 = tmp_io_select;
  assign tmp_tmp_io_select_1 = {2'd0, tmp_tmp_io_select_1_1};
  assign tmp_tmp_weights_ready_1_1 = tmp_weights_ready;
  assign tmp_tmp_weights_ready_1 = {4'd0, tmp_tmp_weights_ready_1_1};
  assign tmp_tmp_weightsAdapted_payload_0_0_0_0 = (tmp_weightsAdapted_payload_0_0_0_0 >>> 128);
  assign tmp_tmp_funcTable_ready_1_1 = tmp_funcTable_ready;
  assign tmp_tmp_funcTable_ready_1 = {3'd0, tmp_tmp_funcTable_ready_1_1};
  StreamFifoHighPerf_2 weightFifo_0 (
    .push_valid               (streamDemux_2_io_outputs_0_valid                  ), //i
    .push_ready               (weightFifo_0_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_0_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_0_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_0_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_0_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_0_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_0_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_0_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_0_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_0_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_0_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_0_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_0_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_0_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_0_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_0_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_0_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_0_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_0_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_0_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_0_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_0_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_0_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_0_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_0_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_0_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_0_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_0_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_0_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_0_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_0_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_0_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_0_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_0_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_0_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_0_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_0_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_0_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_0_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_0_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_0_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_0_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_0_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_0_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_0_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_0_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_0_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_0_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_0_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_0_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_0_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_0_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_0_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_0_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_0_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_0_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_0_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_0_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_0_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_0_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_0_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_0_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_0_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_0_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_0_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_0_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_0_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_0_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_0_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_0_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_0_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_0_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_0_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_0_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_0_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_0_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_0_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_0_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_0_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_0_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_0_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_0_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_0_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_0_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_0_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_0_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_0_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_0_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_0_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_0_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_0_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_0_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_0_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_0_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_0_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_0_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_0_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_0_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_0_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_0_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_0_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_0_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_0_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_0_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_0_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_0_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_0_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_0_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_0_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_0_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_0_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_0_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_0_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_0_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_0_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_0_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_0_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_0_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_0_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_0_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_0_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_0_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_0_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_0_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_0_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_0_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_0_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_0_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_0_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_0_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_0_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_0_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_0_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_0_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_0_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_0_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_0_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_0_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_0_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_0_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_0_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_0_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_0_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_0_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_0_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_0_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_0_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_0_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_0_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_0_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_0_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_0_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_0_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_0_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_0_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_0_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_0_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_0_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_0_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_0_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_0_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_0_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_0_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_0_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_0_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_0_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_0_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_0_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_0_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_0_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_0_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_0_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_0_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_0_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_0_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_0_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_0_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_0_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_0_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_0_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_0_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_0_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_0_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_0_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_0_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_0_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_0_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_0_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_0_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_0_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_0_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_0_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_0_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_0_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_0_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_0_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_0_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_0_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_0_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_0_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_0_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_0_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_0_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_0_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_0_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_0_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_0_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_0_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_0_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_0_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_0_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_0_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_0_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_0_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_0_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_0_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_0_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_0_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_0_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_0_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_0_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_0_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_0_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_0_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_0_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_0_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_0_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_0_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_0_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_0_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_0_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_0_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_0_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_0_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_0_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_0_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_0_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_0_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_0_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_0_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_0_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_0_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_0_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_0_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_0_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_0_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_0_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_0_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_0_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_0_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_0_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_0_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_0_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_0_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_0_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_0_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_0_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_0_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_0_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_0_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_0_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_0_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_0_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_0_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_0_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_0_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_0_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_0_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_0_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_0_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_0_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_0_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_0_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_0_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_0_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_0_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_0_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_0_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_0_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_0_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_0_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_0_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_0_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_0_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_0_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_0_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_0_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_0_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_0_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_0_pop_valid                            ), //o
    .pop_ready                (unit_0_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_0_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_0_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_0_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_0_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_0_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_0_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_0_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_0_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_0_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_0_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_0_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_0_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_0_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_0_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_0_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_0_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_0_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_0_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_0_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_0_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_0_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_0_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_0_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_0_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_0_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_0_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_0_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_0_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_0_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_0_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_0_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_0_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_0_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_0_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_0_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_0_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_0_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_0_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_0_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_0_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_0_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_0_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_0_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_0_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_0_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_0_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_0_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_0_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_0_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_0_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_0_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_0_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_0_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_0_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_0_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_0_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_0_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_0_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_0_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_0_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_0_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_0_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_0_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_0_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_0_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_0_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_0_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_0_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_0_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_0_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_0_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_0_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_0_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_0_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_0_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_0_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_0_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_0_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_0_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_0_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_0_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_0_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_0_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_0_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_0_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_0_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_0_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_0_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_0_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_0_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_0_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_0_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_0_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_0_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_0_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_0_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_0_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_0_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_0_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_0_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_0_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_0_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_0_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_0_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_0_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_0_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_0_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_0_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_0_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_0_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_0_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_0_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_0_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_0_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_0_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_0_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_0_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_0_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_0_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_0_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_0_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_0_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_0_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_0_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_0_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_0_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_0_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_0_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_0_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_0_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_0_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_0_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_0_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_0_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_0_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_0_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_0_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_0_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_0_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_0_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_0_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_0_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_0_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_0_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_0_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_0_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_0_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_0_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_0_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_0_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_0_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_0_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_0_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_0_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_0_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_0_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_0_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_0_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_0_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_0_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_0_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_0_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_0_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_0_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_0_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_0_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_0_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_0_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_0_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_0_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_0_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_0_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_0_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_0_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_0_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_0_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_0_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_0_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_0_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_0_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_0_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_0_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_0_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_0_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_0_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_0_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_0_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_0_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_0_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_0_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_0_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_0_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_0_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_0_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_0_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_0_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_0_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_0_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_0_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_0_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_0_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_0_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_0_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_0_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_0_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_0_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_0_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_0_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_0_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_0_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_0_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_0_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_0_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_0_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_0_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_0_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_0_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_0_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_0_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_0_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_0_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_0_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_0_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_0_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_0_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_0_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_0_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_0_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_0_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_0_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_0_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_0_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_0_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_0_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_0_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_0_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_0_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_0_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_0_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_0_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_0_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_0_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_0_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_0_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_0_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_0_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_0_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_0_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_0_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_0_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_0_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_0_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_0_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_0_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_0_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_0_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_0_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_0_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_0_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_0_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_0_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_0_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_0_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_0_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_0_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_0_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_0_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_0_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_0_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_0_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_0_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_0_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_0_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_0_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_0_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_0_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_0_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_0_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_0_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_0_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_0_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_0_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_0_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_0_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_0_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_0_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_0_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_0_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_1 (
    .push_valid               (streamDemux_2_io_outputs_1_valid                  ), //i
    .push_ready               (weightFifo_1_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_1_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_1_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_1_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_1_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_1_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_1_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_1_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_1_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_1_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_1_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_1_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_1_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_1_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_1_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_1_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_1_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_1_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_1_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_1_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_1_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_1_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_1_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_1_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_1_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_1_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_1_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_1_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_1_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_1_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_1_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_1_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_1_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_1_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_1_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_1_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_1_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_1_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_1_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_1_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_1_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_1_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_1_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_1_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_1_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_1_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_1_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_1_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_1_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_1_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_1_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_1_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_1_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_1_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_1_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_1_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_1_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_1_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_1_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_1_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_1_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_1_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_1_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_1_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_1_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_1_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_1_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_1_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_1_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_1_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_1_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_1_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_1_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_1_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_1_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_1_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_1_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_1_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_1_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_1_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_1_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_1_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_1_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_1_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_1_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_1_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_1_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_1_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_1_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_1_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_1_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_1_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_1_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_1_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_1_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_1_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_1_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_1_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_1_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_1_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_1_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_1_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_1_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_1_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_1_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_1_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_1_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_1_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_1_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_1_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_1_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_1_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_1_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_1_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_1_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_1_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_1_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_1_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_1_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_1_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_1_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_1_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_1_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_1_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_1_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_1_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_1_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_1_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_1_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_1_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_1_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_1_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_1_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_1_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_1_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_1_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_1_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_1_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_1_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_1_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_1_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_1_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_1_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_1_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_1_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_1_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_1_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_1_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_1_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_1_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_1_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_1_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_1_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_1_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_1_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_1_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_1_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_1_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_1_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_1_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_1_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_1_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_1_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_1_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_1_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_1_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_1_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_1_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_1_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_1_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_1_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_1_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_1_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_1_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_1_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_1_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_1_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_1_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_1_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_1_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_1_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_1_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_1_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_1_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_1_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_1_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_1_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_1_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_1_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_1_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_1_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_1_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_1_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_1_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_1_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_1_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_1_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_1_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_1_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_1_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_1_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_1_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_1_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_1_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_1_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_1_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_1_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_1_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_1_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_1_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_1_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_1_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_1_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_1_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_1_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_1_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_1_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_1_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_1_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_1_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_1_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_1_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_1_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_1_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_1_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_1_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_1_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_1_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_1_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_1_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_1_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_1_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_1_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_1_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_1_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_1_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_1_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_1_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_1_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_1_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_1_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_1_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_1_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_1_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_1_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_1_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_1_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_1_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_1_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_1_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_1_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_1_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_1_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_1_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_1_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_1_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_1_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_1_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_1_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_1_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_1_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_1_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_1_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_1_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_1_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_1_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_1_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_1_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_1_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_1_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_1_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_1_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_1_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_1_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_1_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_1_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_1_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_1_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_1_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_1_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_1_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_1_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_1_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_1_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_1_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_1_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_1_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_1_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_1_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_1_pop_valid                            ), //o
    .pop_ready                (unit_1_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_1_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_1_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_1_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_1_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_1_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_1_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_1_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_1_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_1_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_1_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_1_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_1_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_1_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_1_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_1_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_1_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_1_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_1_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_1_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_1_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_1_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_1_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_1_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_1_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_1_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_1_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_1_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_1_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_1_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_1_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_1_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_1_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_1_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_1_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_1_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_1_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_1_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_1_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_1_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_1_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_1_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_1_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_1_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_1_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_1_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_1_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_1_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_1_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_1_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_1_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_1_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_1_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_1_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_1_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_1_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_1_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_1_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_1_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_1_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_1_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_1_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_1_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_1_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_1_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_1_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_1_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_1_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_1_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_1_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_1_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_1_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_1_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_1_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_1_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_1_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_1_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_1_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_1_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_1_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_1_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_1_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_1_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_1_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_1_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_1_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_1_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_1_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_1_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_1_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_1_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_1_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_1_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_1_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_1_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_1_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_1_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_1_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_1_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_1_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_1_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_1_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_1_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_1_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_1_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_1_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_1_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_1_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_1_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_1_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_1_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_1_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_1_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_1_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_1_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_1_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_1_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_1_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_1_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_1_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_1_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_1_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_1_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_1_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_1_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_1_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_1_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_1_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_1_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_1_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_1_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_1_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_1_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_1_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_1_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_1_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_1_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_1_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_1_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_1_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_1_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_1_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_1_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_1_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_1_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_1_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_1_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_1_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_1_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_1_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_1_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_1_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_1_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_1_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_1_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_1_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_1_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_1_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_1_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_1_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_1_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_1_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_1_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_1_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_1_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_1_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_1_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_1_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_1_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_1_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_1_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_1_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_1_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_1_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_1_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_1_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_1_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_1_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_1_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_1_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_1_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_1_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_1_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_1_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_1_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_1_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_1_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_1_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_1_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_1_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_1_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_1_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_1_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_1_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_1_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_1_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_1_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_1_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_1_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_1_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_1_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_1_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_1_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_1_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_1_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_1_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_1_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_1_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_1_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_1_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_1_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_1_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_1_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_1_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_1_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_1_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_1_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_1_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_1_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_1_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_1_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_1_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_1_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_1_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_1_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_1_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_1_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_1_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_1_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_1_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_1_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_1_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_1_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_1_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_1_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_1_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_1_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_1_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_1_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_1_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_1_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_1_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_1_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_1_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_1_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_1_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_1_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_1_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_1_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_1_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_1_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_1_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_1_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_1_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_1_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_1_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_1_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_1_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_1_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_1_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_1_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_1_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_1_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_1_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_1_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_1_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_1_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_1_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_1_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_1_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_1_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_1_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_1_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_1_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_1_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_1_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_1_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_1_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_1_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_1_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_1_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_1_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_1_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_1_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_1_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_1_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_1_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_1_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_1_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_2 (
    .push_valid               (streamDemux_2_io_outputs_2_valid                  ), //i
    .push_ready               (weightFifo_2_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_2_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_2_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_2_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_2_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_2_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_2_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_2_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_2_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_2_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_2_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_2_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_2_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_2_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_2_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_2_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_2_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_2_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_2_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_2_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_2_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_2_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_2_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_2_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_2_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_2_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_2_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_2_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_2_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_2_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_2_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_2_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_2_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_2_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_2_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_2_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_2_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_2_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_2_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_2_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_2_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_2_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_2_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_2_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_2_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_2_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_2_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_2_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_2_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_2_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_2_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_2_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_2_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_2_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_2_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_2_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_2_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_2_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_2_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_2_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_2_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_2_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_2_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_2_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_2_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_2_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_2_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_2_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_2_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_2_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_2_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_2_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_2_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_2_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_2_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_2_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_2_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_2_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_2_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_2_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_2_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_2_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_2_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_2_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_2_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_2_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_2_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_2_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_2_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_2_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_2_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_2_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_2_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_2_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_2_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_2_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_2_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_2_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_2_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_2_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_2_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_2_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_2_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_2_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_2_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_2_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_2_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_2_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_2_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_2_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_2_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_2_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_2_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_2_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_2_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_2_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_2_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_2_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_2_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_2_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_2_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_2_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_2_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_2_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_2_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_2_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_2_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_2_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_2_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_2_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_2_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_2_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_2_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_2_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_2_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_2_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_2_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_2_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_2_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_2_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_2_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_2_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_2_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_2_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_2_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_2_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_2_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_2_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_2_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_2_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_2_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_2_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_2_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_2_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_2_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_2_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_2_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_2_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_2_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_2_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_2_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_2_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_2_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_2_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_2_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_2_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_2_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_2_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_2_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_2_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_2_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_2_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_2_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_2_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_2_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_2_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_2_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_2_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_2_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_2_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_2_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_2_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_2_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_2_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_2_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_2_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_2_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_2_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_2_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_2_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_2_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_2_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_2_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_2_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_2_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_2_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_2_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_2_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_2_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_2_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_2_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_2_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_2_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_2_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_2_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_2_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_2_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_2_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_2_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_2_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_2_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_2_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_2_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_2_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_2_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_2_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_2_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_2_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_2_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_2_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_2_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_2_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_2_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_2_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_2_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_2_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_2_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_2_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_2_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_2_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_2_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_2_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_2_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_2_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_2_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_2_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_2_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_2_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_2_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_2_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_2_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_2_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_2_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_2_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_2_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_2_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_2_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_2_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_2_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_2_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_2_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_2_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_2_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_2_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_2_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_2_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_2_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_2_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_2_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_2_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_2_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_2_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_2_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_2_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_2_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_2_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_2_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_2_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_2_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_2_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_2_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_2_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_2_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_2_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_2_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_2_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_2_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_2_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_2_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_2_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_2_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_2_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_2_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_2_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_2_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_2_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_2_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_2_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_2_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_2_pop_valid                            ), //o
    .pop_ready                (unit_2_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_2_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_2_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_2_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_2_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_2_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_2_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_2_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_2_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_2_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_2_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_2_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_2_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_2_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_2_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_2_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_2_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_2_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_2_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_2_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_2_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_2_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_2_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_2_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_2_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_2_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_2_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_2_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_2_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_2_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_2_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_2_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_2_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_2_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_2_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_2_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_2_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_2_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_2_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_2_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_2_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_2_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_2_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_2_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_2_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_2_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_2_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_2_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_2_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_2_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_2_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_2_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_2_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_2_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_2_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_2_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_2_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_2_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_2_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_2_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_2_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_2_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_2_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_2_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_2_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_2_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_2_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_2_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_2_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_2_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_2_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_2_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_2_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_2_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_2_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_2_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_2_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_2_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_2_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_2_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_2_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_2_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_2_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_2_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_2_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_2_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_2_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_2_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_2_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_2_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_2_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_2_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_2_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_2_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_2_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_2_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_2_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_2_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_2_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_2_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_2_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_2_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_2_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_2_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_2_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_2_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_2_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_2_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_2_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_2_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_2_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_2_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_2_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_2_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_2_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_2_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_2_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_2_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_2_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_2_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_2_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_2_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_2_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_2_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_2_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_2_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_2_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_2_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_2_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_2_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_2_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_2_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_2_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_2_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_2_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_2_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_2_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_2_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_2_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_2_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_2_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_2_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_2_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_2_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_2_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_2_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_2_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_2_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_2_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_2_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_2_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_2_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_2_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_2_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_2_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_2_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_2_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_2_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_2_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_2_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_2_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_2_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_2_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_2_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_2_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_2_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_2_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_2_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_2_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_2_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_2_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_2_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_2_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_2_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_2_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_2_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_2_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_2_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_2_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_2_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_2_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_2_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_2_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_2_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_2_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_2_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_2_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_2_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_2_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_2_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_2_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_2_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_2_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_2_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_2_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_2_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_2_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_2_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_2_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_2_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_2_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_2_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_2_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_2_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_2_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_2_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_2_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_2_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_2_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_2_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_2_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_2_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_2_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_2_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_2_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_2_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_2_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_2_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_2_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_2_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_2_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_2_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_2_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_2_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_2_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_2_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_2_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_2_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_2_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_2_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_2_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_2_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_2_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_2_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_2_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_2_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_2_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_2_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_2_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_2_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_2_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_2_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_2_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_2_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_2_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_2_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_2_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_2_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_2_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_2_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_2_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_2_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_2_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_2_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_2_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_2_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_2_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_2_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_2_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_2_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_2_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_2_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_2_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_2_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_2_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_2_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_2_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_2_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_2_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_2_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_2_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_2_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_2_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_2_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_2_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_2_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_2_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_2_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_2_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_2_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_2_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_2_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_2_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_2_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_2_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_2_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_2_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_2_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_2_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_3 (
    .push_valid               (streamDemux_2_io_outputs_3_valid                  ), //i
    .push_ready               (weightFifo_3_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_3_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_3_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_3_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_3_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_3_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_3_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_3_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_3_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_3_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_3_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_3_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_3_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_3_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_3_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_3_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_3_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_3_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_3_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_3_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_3_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_3_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_3_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_3_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_3_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_3_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_3_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_3_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_3_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_3_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_3_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_3_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_3_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_3_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_3_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_3_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_3_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_3_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_3_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_3_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_3_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_3_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_3_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_3_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_3_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_3_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_3_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_3_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_3_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_3_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_3_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_3_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_3_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_3_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_3_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_3_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_3_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_3_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_3_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_3_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_3_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_3_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_3_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_3_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_3_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_3_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_3_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_3_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_3_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_3_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_3_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_3_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_3_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_3_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_3_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_3_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_3_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_3_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_3_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_3_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_3_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_3_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_3_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_3_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_3_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_3_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_3_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_3_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_3_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_3_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_3_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_3_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_3_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_3_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_3_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_3_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_3_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_3_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_3_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_3_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_3_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_3_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_3_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_3_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_3_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_3_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_3_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_3_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_3_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_3_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_3_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_3_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_3_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_3_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_3_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_3_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_3_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_3_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_3_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_3_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_3_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_3_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_3_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_3_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_3_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_3_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_3_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_3_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_3_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_3_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_3_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_3_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_3_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_3_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_3_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_3_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_3_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_3_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_3_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_3_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_3_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_3_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_3_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_3_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_3_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_3_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_3_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_3_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_3_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_3_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_3_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_3_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_3_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_3_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_3_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_3_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_3_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_3_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_3_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_3_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_3_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_3_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_3_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_3_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_3_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_3_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_3_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_3_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_3_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_3_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_3_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_3_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_3_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_3_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_3_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_3_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_3_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_3_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_3_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_3_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_3_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_3_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_3_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_3_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_3_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_3_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_3_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_3_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_3_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_3_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_3_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_3_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_3_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_3_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_3_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_3_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_3_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_3_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_3_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_3_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_3_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_3_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_3_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_3_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_3_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_3_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_3_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_3_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_3_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_3_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_3_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_3_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_3_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_3_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_3_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_3_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_3_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_3_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_3_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_3_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_3_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_3_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_3_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_3_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_3_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_3_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_3_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_3_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_3_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_3_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_3_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_3_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_3_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_3_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_3_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_3_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_3_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_3_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_3_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_3_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_3_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_3_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_3_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_3_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_3_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_3_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_3_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_3_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_3_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_3_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_3_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_3_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_3_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_3_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_3_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_3_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_3_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_3_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_3_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_3_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_3_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_3_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_3_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_3_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_3_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_3_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_3_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_3_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_3_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_3_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_3_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_3_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_3_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_3_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_3_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_3_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_3_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_3_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_3_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_3_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_3_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_3_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_3_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_3_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_3_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_3_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_3_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_3_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_3_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_3_pop_valid                            ), //o
    .pop_ready                (unit_3_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_3_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_3_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_3_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_3_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_3_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_3_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_3_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_3_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_3_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_3_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_3_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_3_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_3_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_3_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_3_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_3_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_3_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_3_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_3_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_3_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_3_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_3_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_3_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_3_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_3_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_3_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_3_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_3_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_3_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_3_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_3_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_3_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_3_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_3_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_3_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_3_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_3_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_3_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_3_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_3_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_3_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_3_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_3_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_3_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_3_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_3_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_3_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_3_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_3_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_3_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_3_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_3_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_3_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_3_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_3_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_3_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_3_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_3_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_3_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_3_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_3_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_3_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_3_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_3_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_3_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_3_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_3_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_3_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_3_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_3_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_3_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_3_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_3_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_3_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_3_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_3_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_3_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_3_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_3_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_3_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_3_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_3_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_3_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_3_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_3_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_3_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_3_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_3_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_3_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_3_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_3_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_3_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_3_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_3_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_3_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_3_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_3_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_3_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_3_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_3_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_3_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_3_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_3_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_3_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_3_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_3_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_3_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_3_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_3_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_3_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_3_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_3_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_3_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_3_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_3_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_3_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_3_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_3_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_3_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_3_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_3_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_3_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_3_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_3_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_3_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_3_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_3_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_3_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_3_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_3_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_3_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_3_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_3_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_3_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_3_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_3_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_3_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_3_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_3_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_3_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_3_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_3_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_3_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_3_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_3_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_3_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_3_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_3_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_3_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_3_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_3_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_3_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_3_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_3_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_3_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_3_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_3_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_3_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_3_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_3_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_3_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_3_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_3_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_3_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_3_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_3_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_3_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_3_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_3_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_3_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_3_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_3_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_3_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_3_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_3_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_3_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_3_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_3_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_3_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_3_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_3_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_3_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_3_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_3_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_3_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_3_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_3_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_3_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_3_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_3_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_3_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_3_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_3_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_3_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_3_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_3_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_3_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_3_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_3_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_3_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_3_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_3_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_3_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_3_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_3_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_3_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_3_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_3_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_3_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_3_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_3_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_3_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_3_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_3_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_3_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_3_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_3_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_3_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_3_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_3_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_3_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_3_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_3_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_3_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_3_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_3_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_3_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_3_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_3_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_3_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_3_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_3_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_3_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_3_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_3_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_3_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_3_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_3_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_3_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_3_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_3_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_3_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_3_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_3_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_3_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_3_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_3_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_3_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_3_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_3_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_3_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_3_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_3_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_3_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_3_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_3_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_3_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_3_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_3_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_3_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_3_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_3_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_3_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_3_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_3_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_3_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_3_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_3_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_3_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_3_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_3_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_3_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_3_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_3_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_3_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_3_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_3_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_3_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_3_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_3_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_3_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_3_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_3_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_3_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_3_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_3_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_3_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_3_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_4 (
    .push_valid               (streamDemux_2_io_outputs_4_valid                  ), //i
    .push_ready               (weightFifo_4_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_4_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_4_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_4_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_4_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_4_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_4_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_4_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_4_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_4_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_4_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_4_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_4_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_4_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_4_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_4_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_4_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_4_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_4_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_4_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_4_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_4_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_4_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_4_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_4_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_4_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_4_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_4_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_4_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_4_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_4_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_4_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_4_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_4_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_4_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_4_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_4_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_4_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_4_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_4_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_4_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_4_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_4_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_4_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_4_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_4_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_4_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_4_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_4_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_4_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_4_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_4_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_4_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_4_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_4_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_4_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_4_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_4_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_4_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_4_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_4_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_4_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_4_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_4_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_4_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_4_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_4_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_4_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_4_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_4_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_4_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_4_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_4_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_4_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_4_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_4_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_4_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_4_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_4_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_4_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_4_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_4_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_4_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_4_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_4_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_4_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_4_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_4_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_4_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_4_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_4_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_4_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_4_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_4_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_4_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_4_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_4_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_4_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_4_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_4_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_4_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_4_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_4_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_4_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_4_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_4_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_4_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_4_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_4_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_4_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_4_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_4_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_4_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_4_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_4_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_4_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_4_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_4_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_4_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_4_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_4_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_4_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_4_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_4_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_4_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_4_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_4_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_4_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_4_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_4_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_4_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_4_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_4_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_4_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_4_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_4_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_4_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_4_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_4_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_4_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_4_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_4_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_4_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_4_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_4_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_4_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_4_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_4_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_4_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_4_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_4_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_4_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_4_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_4_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_4_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_4_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_4_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_4_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_4_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_4_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_4_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_4_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_4_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_4_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_4_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_4_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_4_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_4_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_4_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_4_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_4_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_4_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_4_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_4_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_4_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_4_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_4_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_4_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_4_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_4_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_4_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_4_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_4_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_4_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_4_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_4_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_4_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_4_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_4_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_4_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_4_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_4_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_4_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_4_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_4_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_4_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_4_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_4_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_4_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_4_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_4_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_4_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_4_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_4_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_4_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_4_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_4_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_4_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_4_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_4_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_4_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_4_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_4_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_4_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_4_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_4_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_4_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_4_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_4_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_4_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_4_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_4_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_4_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_4_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_4_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_4_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_4_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_4_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_4_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_4_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_4_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_4_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_4_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_4_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_4_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_4_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_4_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_4_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_4_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_4_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_4_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_4_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_4_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_4_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_4_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_4_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_4_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_4_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_4_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_4_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_4_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_4_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_4_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_4_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_4_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_4_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_4_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_4_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_4_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_4_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_4_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_4_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_4_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_4_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_4_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_4_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_4_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_4_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_4_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_4_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_4_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_4_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_4_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_4_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_4_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_4_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_4_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_4_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_4_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_4_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_4_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_4_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_4_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_4_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_4_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_4_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_4_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_4_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_4_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_4_pop_valid                            ), //o
    .pop_ready                (unit_4_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_4_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_4_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_4_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_4_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_4_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_4_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_4_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_4_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_4_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_4_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_4_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_4_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_4_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_4_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_4_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_4_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_4_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_4_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_4_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_4_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_4_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_4_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_4_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_4_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_4_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_4_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_4_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_4_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_4_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_4_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_4_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_4_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_4_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_4_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_4_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_4_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_4_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_4_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_4_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_4_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_4_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_4_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_4_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_4_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_4_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_4_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_4_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_4_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_4_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_4_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_4_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_4_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_4_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_4_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_4_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_4_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_4_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_4_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_4_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_4_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_4_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_4_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_4_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_4_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_4_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_4_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_4_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_4_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_4_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_4_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_4_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_4_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_4_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_4_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_4_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_4_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_4_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_4_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_4_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_4_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_4_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_4_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_4_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_4_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_4_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_4_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_4_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_4_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_4_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_4_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_4_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_4_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_4_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_4_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_4_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_4_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_4_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_4_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_4_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_4_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_4_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_4_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_4_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_4_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_4_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_4_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_4_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_4_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_4_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_4_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_4_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_4_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_4_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_4_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_4_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_4_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_4_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_4_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_4_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_4_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_4_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_4_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_4_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_4_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_4_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_4_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_4_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_4_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_4_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_4_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_4_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_4_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_4_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_4_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_4_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_4_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_4_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_4_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_4_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_4_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_4_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_4_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_4_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_4_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_4_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_4_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_4_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_4_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_4_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_4_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_4_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_4_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_4_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_4_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_4_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_4_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_4_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_4_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_4_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_4_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_4_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_4_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_4_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_4_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_4_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_4_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_4_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_4_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_4_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_4_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_4_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_4_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_4_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_4_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_4_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_4_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_4_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_4_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_4_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_4_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_4_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_4_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_4_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_4_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_4_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_4_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_4_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_4_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_4_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_4_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_4_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_4_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_4_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_4_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_4_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_4_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_4_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_4_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_4_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_4_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_4_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_4_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_4_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_4_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_4_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_4_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_4_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_4_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_4_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_4_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_4_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_4_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_4_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_4_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_4_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_4_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_4_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_4_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_4_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_4_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_4_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_4_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_4_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_4_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_4_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_4_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_4_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_4_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_4_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_4_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_4_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_4_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_4_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_4_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_4_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_4_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_4_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_4_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_4_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_4_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_4_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_4_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_4_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_4_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_4_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_4_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_4_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_4_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_4_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_4_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_4_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_4_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_4_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_4_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_4_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_4_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_4_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_4_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_4_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_4_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_4_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_4_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_4_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_4_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_4_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_4_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_4_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_4_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_4_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_4_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_4_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_4_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_4_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_4_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_4_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_4_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_4_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_4_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_4_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_4_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_4_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_4_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_4_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_4_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_4_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_4_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_4_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_4_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_5 (
    .push_valid               (streamDemux_2_io_outputs_5_valid                  ), //i
    .push_ready               (weightFifo_5_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_5_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_5_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_5_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_5_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_5_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_5_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_5_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_5_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_5_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_5_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_5_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_5_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_5_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_5_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_5_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_5_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_5_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_5_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_5_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_5_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_5_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_5_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_5_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_5_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_5_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_5_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_5_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_5_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_5_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_5_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_5_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_5_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_5_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_5_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_5_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_5_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_5_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_5_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_5_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_5_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_5_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_5_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_5_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_5_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_5_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_5_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_5_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_5_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_5_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_5_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_5_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_5_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_5_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_5_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_5_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_5_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_5_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_5_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_5_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_5_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_5_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_5_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_5_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_5_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_5_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_5_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_5_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_5_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_5_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_5_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_5_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_5_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_5_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_5_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_5_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_5_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_5_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_5_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_5_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_5_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_5_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_5_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_5_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_5_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_5_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_5_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_5_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_5_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_5_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_5_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_5_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_5_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_5_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_5_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_5_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_5_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_5_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_5_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_5_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_5_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_5_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_5_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_5_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_5_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_5_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_5_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_5_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_5_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_5_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_5_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_5_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_5_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_5_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_5_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_5_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_5_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_5_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_5_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_5_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_5_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_5_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_5_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_5_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_5_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_5_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_5_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_5_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_5_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_5_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_5_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_5_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_5_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_5_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_5_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_5_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_5_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_5_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_5_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_5_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_5_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_5_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_5_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_5_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_5_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_5_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_5_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_5_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_5_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_5_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_5_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_5_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_5_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_5_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_5_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_5_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_5_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_5_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_5_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_5_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_5_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_5_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_5_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_5_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_5_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_5_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_5_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_5_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_5_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_5_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_5_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_5_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_5_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_5_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_5_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_5_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_5_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_5_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_5_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_5_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_5_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_5_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_5_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_5_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_5_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_5_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_5_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_5_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_5_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_5_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_5_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_5_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_5_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_5_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_5_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_5_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_5_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_5_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_5_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_5_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_5_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_5_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_5_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_5_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_5_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_5_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_5_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_5_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_5_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_5_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_5_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_5_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_5_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_5_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_5_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_5_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_5_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_5_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_5_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_5_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_5_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_5_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_5_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_5_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_5_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_5_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_5_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_5_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_5_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_5_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_5_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_5_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_5_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_5_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_5_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_5_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_5_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_5_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_5_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_5_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_5_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_5_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_5_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_5_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_5_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_5_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_5_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_5_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_5_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_5_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_5_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_5_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_5_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_5_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_5_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_5_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_5_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_5_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_5_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_5_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_5_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_5_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_5_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_5_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_5_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_5_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_5_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_5_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_5_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_5_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_5_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_5_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_5_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_5_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_5_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_5_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_5_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_5_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_5_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_5_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_5_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_5_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_5_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_5_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_5_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_5_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_5_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_5_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_5_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_5_pop_valid                            ), //o
    .pop_ready                (unit_5_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_5_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_5_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_5_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_5_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_5_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_5_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_5_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_5_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_5_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_5_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_5_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_5_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_5_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_5_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_5_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_5_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_5_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_5_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_5_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_5_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_5_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_5_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_5_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_5_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_5_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_5_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_5_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_5_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_5_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_5_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_5_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_5_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_5_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_5_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_5_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_5_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_5_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_5_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_5_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_5_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_5_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_5_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_5_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_5_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_5_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_5_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_5_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_5_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_5_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_5_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_5_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_5_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_5_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_5_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_5_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_5_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_5_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_5_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_5_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_5_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_5_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_5_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_5_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_5_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_5_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_5_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_5_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_5_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_5_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_5_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_5_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_5_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_5_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_5_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_5_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_5_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_5_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_5_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_5_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_5_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_5_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_5_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_5_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_5_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_5_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_5_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_5_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_5_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_5_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_5_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_5_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_5_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_5_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_5_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_5_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_5_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_5_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_5_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_5_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_5_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_5_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_5_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_5_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_5_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_5_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_5_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_5_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_5_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_5_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_5_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_5_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_5_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_5_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_5_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_5_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_5_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_5_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_5_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_5_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_5_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_5_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_5_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_5_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_5_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_5_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_5_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_5_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_5_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_5_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_5_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_5_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_5_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_5_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_5_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_5_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_5_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_5_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_5_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_5_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_5_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_5_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_5_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_5_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_5_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_5_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_5_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_5_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_5_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_5_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_5_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_5_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_5_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_5_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_5_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_5_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_5_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_5_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_5_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_5_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_5_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_5_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_5_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_5_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_5_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_5_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_5_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_5_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_5_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_5_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_5_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_5_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_5_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_5_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_5_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_5_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_5_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_5_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_5_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_5_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_5_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_5_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_5_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_5_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_5_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_5_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_5_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_5_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_5_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_5_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_5_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_5_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_5_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_5_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_5_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_5_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_5_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_5_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_5_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_5_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_5_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_5_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_5_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_5_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_5_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_5_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_5_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_5_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_5_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_5_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_5_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_5_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_5_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_5_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_5_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_5_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_5_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_5_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_5_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_5_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_5_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_5_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_5_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_5_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_5_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_5_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_5_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_5_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_5_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_5_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_5_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_5_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_5_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_5_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_5_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_5_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_5_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_5_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_5_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_5_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_5_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_5_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_5_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_5_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_5_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_5_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_5_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_5_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_5_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_5_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_5_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_5_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_5_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_5_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_5_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_5_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_5_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_5_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_5_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_5_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_5_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_5_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_5_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_5_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_5_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_5_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_5_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_5_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_5_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_5_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_5_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_5_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_5_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_5_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_5_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_5_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_5_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_5_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_5_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_5_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_5_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_5_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_5_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_5_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_5_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_5_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_5_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_5_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_5_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_6 (
    .push_valid               (streamDemux_2_io_outputs_6_valid                  ), //i
    .push_ready               (weightFifo_6_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_6_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_6_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_6_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_6_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_6_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_6_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_6_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_6_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_6_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_6_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_6_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_6_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_6_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_6_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_6_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_6_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_6_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_6_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_6_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_6_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_6_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_6_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_6_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_6_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_6_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_6_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_6_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_6_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_6_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_6_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_6_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_6_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_6_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_6_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_6_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_6_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_6_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_6_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_6_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_6_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_6_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_6_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_6_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_6_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_6_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_6_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_6_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_6_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_6_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_6_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_6_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_6_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_6_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_6_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_6_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_6_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_6_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_6_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_6_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_6_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_6_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_6_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_6_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_6_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_6_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_6_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_6_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_6_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_6_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_6_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_6_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_6_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_6_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_6_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_6_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_6_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_6_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_6_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_6_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_6_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_6_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_6_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_6_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_6_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_6_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_6_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_6_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_6_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_6_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_6_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_6_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_6_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_6_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_6_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_6_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_6_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_6_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_6_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_6_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_6_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_6_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_6_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_6_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_6_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_6_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_6_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_6_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_6_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_6_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_6_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_6_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_6_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_6_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_6_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_6_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_6_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_6_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_6_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_6_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_6_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_6_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_6_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_6_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_6_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_6_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_6_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_6_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_6_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_6_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_6_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_6_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_6_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_6_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_6_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_6_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_6_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_6_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_6_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_6_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_6_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_6_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_6_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_6_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_6_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_6_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_6_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_6_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_6_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_6_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_6_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_6_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_6_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_6_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_6_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_6_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_6_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_6_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_6_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_6_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_6_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_6_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_6_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_6_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_6_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_6_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_6_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_6_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_6_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_6_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_6_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_6_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_6_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_6_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_6_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_6_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_6_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_6_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_6_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_6_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_6_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_6_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_6_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_6_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_6_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_6_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_6_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_6_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_6_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_6_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_6_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_6_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_6_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_6_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_6_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_6_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_6_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_6_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_6_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_6_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_6_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_6_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_6_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_6_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_6_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_6_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_6_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_6_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_6_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_6_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_6_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_6_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_6_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_6_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_6_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_6_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_6_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_6_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_6_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_6_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_6_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_6_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_6_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_6_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_6_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_6_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_6_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_6_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_6_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_6_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_6_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_6_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_6_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_6_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_6_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_6_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_6_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_6_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_6_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_6_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_6_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_6_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_6_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_6_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_6_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_6_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_6_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_6_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_6_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_6_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_6_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_6_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_6_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_6_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_6_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_6_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_6_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_6_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_6_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_6_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_6_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_6_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_6_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_6_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_6_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_6_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_6_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_6_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_6_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_6_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_6_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_6_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_6_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_6_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_6_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_6_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_6_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_6_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_6_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_6_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_6_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_6_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_6_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_6_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_6_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_6_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_6_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_6_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_6_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_6_pop_valid                            ), //o
    .pop_ready                (unit_6_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_6_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_6_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_6_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_6_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_6_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_6_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_6_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_6_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_6_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_6_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_6_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_6_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_6_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_6_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_6_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_6_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_6_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_6_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_6_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_6_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_6_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_6_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_6_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_6_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_6_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_6_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_6_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_6_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_6_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_6_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_6_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_6_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_6_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_6_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_6_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_6_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_6_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_6_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_6_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_6_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_6_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_6_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_6_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_6_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_6_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_6_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_6_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_6_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_6_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_6_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_6_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_6_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_6_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_6_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_6_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_6_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_6_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_6_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_6_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_6_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_6_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_6_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_6_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_6_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_6_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_6_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_6_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_6_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_6_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_6_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_6_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_6_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_6_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_6_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_6_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_6_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_6_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_6_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_6_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_6_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_6_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_6_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_6_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_6_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_6_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_6_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_6_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_6_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_6_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_6_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_6_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_6_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_6_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_6_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_6_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_6_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_6_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_6_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_6_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_6_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_6_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_6_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_6_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_6_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_6_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_6_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_6_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_6_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_6_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_6_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_6_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_6_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_6_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_6_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_6_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_6_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_6_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_6_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_6_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_6_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_6_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_6_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_6_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_6_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_6_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_6_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_6_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_6_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_6_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_6_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_6_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_6_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_6_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_6_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_6_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_6_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_6_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_6_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_6_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_6_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_6_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_6_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_6_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_6_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_6_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_6_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_6_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_6_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_6_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_6_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_6_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_6_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_6_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_6_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_6_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_6_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_6_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_6_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_6_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_6_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_6_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_6_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_6_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_6_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_6_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_6_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_6_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_6_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_6_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_6_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_6_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_6_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_6_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_6_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_6_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_6_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_6_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_6_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_6_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_6_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_6_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_6_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_6_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_6_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_6_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_6_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_6_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_6_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_6_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_6_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_6_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_6_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_6_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_6_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_6_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_6_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_6_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_6_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_6_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_6_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_6_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_6_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_6_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_6_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_6_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_6_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_6_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_6_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_6_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_6_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_6_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_6_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_6_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_6_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_6_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_6_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_6_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_6_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_6_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_6_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_6_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_6_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_6_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_6_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_6_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_6_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_6_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_6_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_6_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_6_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_6_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_6_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_6_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_6_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_6_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_6_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_6_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_6_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_6_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_6_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_6_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_6_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_6_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_6_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_6_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_6_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_6_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_6_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_6_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_6_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_6_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_6_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_6_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_6_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_6_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_6_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_6_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_6_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_6_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_6_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_6_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_6_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_6_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_6_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_6_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_6_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_6_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_6_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_6_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_6_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_6_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_6_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_6_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_6_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_6_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_6_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_6_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_6_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_6_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_6_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_6_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_6_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_6_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_6_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_6_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_6_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_6_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_6_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  StreamFifoHighPerf_2 weightFifo_7 (
    .push_valid               (streamDemux_2_io_outputs_7_valid                  ), //i
    .push_ready               (weightFifo_7_push_ready                           ), //o
    .push_payload_0_0_0_0     (streamDemux_2_io_outputs_7_payload_0_0_0_0[7:0]   ), //i
    .push_payload_0_0_0_1     (streamDemux_2_io_outputs_7_payload_0_0_0_1[7:0]   ), //i
    .push_payload_0_0_0_2     (streamDemux_2_io_outputs_7_payload_0_0_0_2[7:0]   ), //i
    .push_payload_0_0_0_3     (streamDemux_2_io_outputs_7_payload_0_0_0_3[7:0]   ), //i
    .push_payload_0_0_0_4     (streamDemux_2_io_outputs_7_payload_0_0_0_4[7:0]   ), //i
    .push_payload_0_0_0_5     (streamDemux_2_io_outputs_7_payload_0_0_0_5[7:0]   ), //i
    .push_payload_0_0_0_6     (streamDemux_2_io_outputs_7_payload_0_0_0_6[7:0]   ), //i
    .push_payload_0_0_0_7     (streamDemux_2_io_outputs_7_payload_0_0_0_7[7:0]   ), //i
    .push_payload_0_0_0_8     (streamDemux_2_io_outputs_7_payload_0_0_0_8[7:0]   ), //i
    .push_payload_0_0_0_9     (streamDemux_2_io_outputs_7_payload_0_0_0_9[7:0]   ), //i
    .push_payload_0_0_0_10    (streamDemux_2_io_outputs_7_payload_0_0_0_10[7:0]  ), //i
    .push_payload_0_0_0_11    (streamDemux_2_io_outputs_7_payload_0_0_0_11[7:0]  ), //i
    .push_payload_0_0_0_12    (streamDemux_2_io_outputs_7_payload_0_0_0_12[7:0]  ), //i
    .push_payload_0_0_0_13    (streamDemux_2_io_outputs_7_payload_0_0_0_13[7:0]  ), //i
    .push_payload_0_0_0_14    (streamDemux_2_io_outputs_7_payload_0_0_0_14[7:0]  ), //i
    .push_payload_0_0_0_15    (streamDemux_2_io_outputs_7_payload_0_0_0_15[7:0]  ), //i
    .push_payload_0_0_1_0     (streamDemux_2_io_outputs_7_payload_0_0_1_0[7:0]   ), //i
    .push_payload_0_0_1_1     (streamDemux_2_io_outputs_7_payload_0_0_1_1[7:0]   ), //i
    .push_payload_0_0_1_2     (streamDemux_2_io_outputs_7_payload_0_0_1_2[7:0]   ), //i
    .push_payload_0_0_1_3     (streamDemux_2_io_outputs_7_payload_0_0_1_3[7:0]   ), //i
    .push_payload_0_0_1_4     (streamDemux_2_io_outputs_7_payload_0_0_1_4[7:0]   ), //i
    .push_payload_0_0_1_5     (streamDemux_2_io_outputs_7_payload_0_0_1_5[7:0]   ), //i
    .push_payload_0_0_1_6     (streamDemux_2_io_outputs_7_payload_0_0_1_6[7:0]   ), //i
    .push_payload_0_0_1_7     (streamDemux_2_io_outputs_7_payload_0_0_1_7[7:0]   ), //i
    .push_payload_0_0_1_8     (streamDemux_2_io_outputs_7_payload_0_0_1_8[7:0]   ), //i
    .push_payload_0_0_1_9     (streamDemux_2_io_outputs_7_payload_0_0_1_9[7:0]   ), //i
    .push_payload_0_0_1_10    (streamDemux_2_io_outputs_7_payload_0_0_1_10[7:0]  ), //i
    .push_payload_0_0_1_11    (streamDemux_2_io_outputs_7_payload_0_0_1_11[7:0]  ), //i
    .push_payload_0_0_1_12    (streamDemux_2_io_outputs_7_payload_0_0_1_12[7:0]  ), //i
    .push_payload_0_0_1_13    (streamDemux_2_io_outputs_7_payload_0_0_1_13[7:0]  ), //i
    .push_payload_0_0_1_14    (streamDemux_2_io_outputs_7_payload_0_0_1_14[7:0]  ), //i
    .push_payload_0_0_1_15    (streamDemux_2_io_outputs_7_payload_0_0_1_15[7:0]  ), //i
    .push_payload_0_0_2_0     (streamDemux_2_io_outputs_7_payload_0_0_2_0[7:0]   ), //i
    .push_payload_0_0_2_1     (streamDemux_2_io_outputs_7_payload_0_0_2_1[7:0]   ), //i
    .push_payload_0_0_2_2     (streamDemux_2_io_outputs_7_payload_0_0_2_2[7:0]   ), //i
    .push_payload_0_0_2_3     (streamDemux_2_io_outputs_7_payload_0_0_2_3[7:0]   ), //i
    .push_payload_0_0_2_4     (streamDemux_2_io_outputs_7_payload_0_0_2_4[7:0]   ), //i
    .push_payload_0_0_2_5     (streamDemux_2_io_outputs_7_payload_0_0_2_5[7:0]   ), //i
    .push_payload_0_0_2_6     (streamDemux_2_io_outputs_7_payload_0_0_2_6[7:0]   ), //i
    .push_payload_0_0_2_7     (streamDemux_2_io_outputs_7_payload_0_0_2_7[7:0]   ), //i
    .push_payload_0_0_2_8     (streamDemux_2_io_outputs_7_payload_0_0_2_8[7:0]   ), //i
    .push_payload_0_0_2_9     (streamDemux_2_io_outputs_7_payload_0_0_2_9[7:0]   ), //i
    .push_payload_0_0_2_10    (streamDemux_2_io_outputs_7_payload_0_0_2_10[7:0]  ), //i
    .push_payload_0_0_2_11    (streamDemux_2_io_outputs_7_payload_0_0_2_11[7:0]  ), //i
    .push_payload_0_0_2_12    (streamDemux_2_io_outputs_7_payload_0_0_2_12[7:0]  ), //i
    .push_payload_0_0_2_13    (streamDemux_2_io_outputs_7_payload_0_0_2_13[7:0]  ), //i
    .push_payload_0_0_2_14    (streamDemux_2_io_outputs_7_payload_0_0_2_14[7:0]  ), //i
    .push_payload_0_0_2_15    (streamDemux_2_io_outputs_7_payload_0_0_2_15[7:0]  ), //i
    .push_payload_0_1_0_0     (streamDemux_2_io_outputs_7_payload_0_1_0_0[7:0]   ), //i
    .push_payload_0_1_0_1     (streamDemux_2_io_outputs_7_payload_0_1_0_1[7:0]   ), //i
    .push_payload_0_1_0_2     (streamDemux_2_io_outputs_7_payload_0_1_0_2[7:0]   ), //i
    .push_payload_0_1_0_3     (streamDemux_2_io_outputs_7_payload_0_1_0_3[7:0]   ), //i
    .push_payload_0_1_0_4     (streamDemux_2_io_outputs_7_payload_0_1_0_4[7:0]   ), //i
    .push_payload_0_1_0_5     (streamDemux_2_io_outputs_7_payload_0_1_0_5[7:0]   ), //i
    .push_payload_0_1_0_6     (streamDemux_2_io_outputs_7_payload_0_1_0_6[7:0]   ), //i
    .push_payload_0_1_0_7     (streamDemux_2_io_outputs_7_payload_0_1_0_7[7:0]   ), //i
    .push_payload_0_1_0_8     (streamDemux_2_io_outputs_7_payload_0_1_0_8[7:0]   ), //i
    .push_payload_0_1_0_9     (streamDemux_2_io_outputs_7_payload_0_1_0_9[7:0]   ), //i
    .push_payload_0_1_0_10    (streamDemux_2_io_outputs_7_payload_0_1_0_10[7:0]  ), //i
    .push_payload_0_1_0_11    (streamDemux_2_io_outputs_7_payload_0_1_0_11[7:0]  ), //i
    .push_payload_0_1_0_12    (streamDemux_2_io_outputs_7_payload_0_1_0_12[7:0]  ), //i
    .push_payload_0_1_0_13    (streamDemux_2_io_outputs_7_payload_0_1_0_13[7:0]  ), //i
    .push_payload_0_1_0_14    (streamDemux_2_io_outputs_7_payload_0_1_0_14[7:0]  ), //i
    .push_payload_0_1_0_15    (streamDemux_2_io_outputs_7_payload_0_1_0_15[7:0]  ), //i
    .push_payload_0_1_1_0     (streamDemux_2_io_outputs_7_payload_0_1_1_0[7:0]   ), //i
    .push_payload_0_1_1_1     (streamDemux_2_io_outputs_7_payload_0_1_1_1[7:0]   ), //i
    .push_payload_0_1_1_2     (streamDemux_2_io_outputs_7_payload_0_1_1_2[7:0]   ), //i
    .push_payload_0_1_1_3     (streamDemux_2_io_outputs_7_payload_0_1_1_3[7:0]   ), //i
    .push_payload_0_1_1_4     (streamDemux_2_io_outputs_7_payload_0_1_1_4[7:0]   ), //i
    .push_payload_0_1_1_5     (streamDemux_2_io_outputs_7_payload_0_1_1_5[7:0]   ), //i
    .push_payload_0_1_1_6     (streamDemux_2_io_outputs_7_payload_0_1_1_6[7:0]   ), //i
    .push_payload_0_1_1_7     (streamDemux_2_io_outputs_7_payload_0_1_1_7[7:0]   ), //i
    .push_payload_0_1_1_8     (streamDemux_2_io_outputs_7_payload_0_1_1_8[7:0]   ), //i
    .push_payload_0_1_1_9     (streamDemux_2_io_outputs_7_payload_0_1_1_9[7:0]   ), //i
    .push_payload_0_1_1_10    (streamDemux_2_io_outputs_7_payload_0_1_1_10[7:0]  ), //i
    .push_payload_0_1_1_11    (streamDemux_2_io_outputs_7_payload_0_1_1_11[7:0]  ), //i
    .push_payload_0_1_1_12    (streamDemux_2_io_outputs_7_payload_0_1_1_12[7:0]  ), //i
    .push_payload_0_1_1_13    (streamDemux_2_io_outputs_7_payload_0_1_1_13[7:0]  ), //i
    .push_payload_0_1_1_14    (streamDemux_2_io_outputs_7_payload_0_1_1_14[7:0]  ), //i
    .push_payload_0_1_1_15    (streamDemux_2_io_outputs_7_payload_0_1_1_15[7:0]  ), //i
    .push_payload_0_1_2_0     (streamDemux_2_io_outputs_7_payload_0_1_2_0[7:0]   ), //i
    .push_payload_0_1_2_1     (streamDemux_2_io_outputs_7_payload_0_1_2_1[7:0]   ), //i
    .push_payload_0_1_2_2     (streamDemux_2_io_outputs_7_payload_0_1_2_2[7:0]   ), //i
    .push_payload_0_1_2_3     (streamDemux_2_io_outputs_7_payload_0_1_2_3[7:0]   ), //i
    .push_payload_0_1_2_4     (streamDemux_2_io_outputs_7_payload_0_1_2_4[7:0]   ), //i
    .push_payload_0_1_2_5     (streamDemux_2_io_outputs_7_payload_0_1_2_5[7:0]   ), //i
    .push_payload_0_1_2_6     (streamDemux_2_io_outputs_7_payload_0_1_2_6[7:0]   ), //i
    .push_payload_0_1_2_7     (streamDemux_2_io_outputs_7_payload_0_1_2_7[7:0]   ), //i
    .push_payload_0_1_2_8     (streamDemux_2_io_outputs_7_payload_0_1_2_8[7:0]   ), //i
    .push_payload_0_1_2_9     (streamDemux_2_io_outputs_7_payload_0_1_2_9[7:0]   ), //i
    .push_payload_0_1_2_10    (streamDemux_2_io_outputs_7_payload_0_1_2_10[7:0]  ), //i
    .push_payload_0_1_2_11    (streamDemux_2_io_outputs_7_payload_0_1_2_11[7:0]  ), //i
    .push_payload_0_1_2_12    (streamDemux_2_io_outputs_7_payload_0_1_2_12[7:0]  ), //i
    .push_payload_0_1_2_13    (streamDemux_2_io_outputs_7_payload_0_1_2_13[7:0]  ), //i
    .push_payload_0_1_2_14    (streamDemux_2_io_outputs_7_payload_0_1_2_14[7:0]  ), //i
    .push_payload_0_1_2_15    (streamDemux_2_io_outputs_7_payload_0_1_2_15[7:0]  ), //i
    .push_payload_0_2_0_0     (streamDemux_2_io_outputs_7_payload_0_2_0_0[7:0]   ), //i
    .push_payload_0_2_0_1     (streamDemux_2_io_outputs_7_payload_0_2_0_1[7:0]   ), //i
    .push_payload_0_2_0_2     (streamDemux_2_io_outputs_7_payload_0_2_0_2[7:0]   ), //i
    .push_payload_0_2_0_3     (streamDemux_2_io_outputs_7_payload_0_2_0_3[7:0]   ), //i
    .push_payload_0_2_0_4     (streamDemux_2_io_outputs_7_payload_0_2_0_4[7:0]   ), //i
    .push_payload_0_2_0_5     (streamDemux_2_io_outputs_7_payload_0_2_0_5[7:0]   ), //i
    .push_payload_0_2_0_6     (streamDemux_2_io_outputs_7_payload_0_2_0_6[7:0]   ), //i
    .push_payload_0_2_0_7     (streamDemux_2_io_outputs_7_payload_0_2_0_7[7:0]   ), //i
    .push_payload_0_2_0_8     (streamDemux_2_io_outputs_7_payload_0_2_0_8[7:0]   ), //i
    .push_payload_0_2_0_9     (streamDemux_2_io_outputs_7_payload_0_2_0_9[7:0]   ), //i
    .push_payload_0_2_0_10    (streamDemux_2_io_outputs_7_payload_0_2_0_10[7:0]  ), //i
    .push_payload_0_2_0_11    (streamDemux_2_io_outputs_7_payload_0_2_0_11[7:0]  ), //i
    .push_payload_0_2_0_12    (streamDemux_2_io_outputs_7_payload_0_2_0_12[7:0]  ), //i
    .push_payload_0_2_0_13    (streamDemux_2_io_outputs_7_payload_0_2_0_13[7:0]  ), //i
    .push_payload_0_2_0_14    (streamDemux_2_io_outputs_7_payload_0_2_0_14[7:0]  ), //i
    .push_payload_0_2_0_15    (streamDemux_2_io_outputs_7_payload_0_2_0_15[7:0]  ), //i
    .push_payload_0_2_1_0     (streamDemux_2_io_outputs_7_payload_0_2_1_0[7:0]   ), //i
    .push_payload_0_2_1_1     (streamDemux_2_io_outputs_7_payload_0_2_1_1[7:0]   ), //i
    .push_payload_0_2_1_2     (streamDemux_2_io_outputs_7_payload_0_2_1_2[7:0]   ), //i
    .push_payload_0_2_1_3     (streamDemux_2_io_outputs_7_payload_0_2_1_3[7:0]   ), //i
    .push_payload_0_2_1_4     (streamDemux_2_io_outputs_7_payload_0_2_1_4[7:0]   ), //i
    .push_payload_0_2_1_5     (streamDemux_2_io_outputs_7_payload_0_2_1_5[7:0]   ), //i
    .push_payload_0_2_1_6     (streamDemux_2_io_outputs_7_payload_0_2_1_6[7:0]   ), //i
    .push_payload_0_2_1_7     (streamDemux_2_io_outputs_7_payload_0_2_1_7[7:0]   ), //i
    .push_payload_0_2_1_8     (streamDemux_2_io_outputs_7_payload_0_2_1_8[7:0]   ), //i
    .push_payload_0_2_1_9     (streamDemux_2_io_outputs_7_payload_0_2_1_9[7:0]   ), //i
    .push_payload_0_2_1_10    (streamDemux_2_io_outputs_7_payload_0_2_1_10[7:0]  ), //i
    .push_payload_0_2_1_11    (streamDemux_2_io_outputs_7_payload_0_2_1_11[7:0]  ), //i
    .push_payload_0_2_1_12    (streamDemux_2_io_outputs_7_payload_0_2_1_12[7:0]  ), //i
    .push_payload_0_2_1_13    (streamDemux_2_io_outputs_7_payload_0_2_1_13[7:0]  ), //i
    .push_payload_0_2_1_14    (streamDemux_2_io_outputs_7_payload_0_2_1_14[7:0]  ), //i
    .push_payload_0_2_1_15    (streamDemux_2_io_outputs_7_payload_0_2_1_15[7:0]  ), //i
    .push_payload_0_2_2_0     (streamDemux_2_io_outputs_7_payload_0_2_2_0[7:0]   ), //i
    .push_payload_0_2_2_1     (streamDemux_2_io_outputs_7_payload_0_2_2_1[7:0]   ), //i
    .push_payload_0_2_2_2     (streamDemux_2_io_outputs_7_payload_0_2_2_2[7:0]   ), //i
    .push_payload_0_2_2_3     (streamDemux_2_io_outputs_7_payload_0_2_2_3[7:0]   ), //i
    .push_payload_0_2_2_4     (streamDemux_2_io_outputs_7_payload_0_2_2_4[7:0]   ), //i
    .push_payload_0_2_2_5     (streamDemux_2_io_outputs_7_payload_0_2_2_5[7:0]   ), //i
    .push_payload_0_2_2_6     (streamDemux_2_io_outputs_7_payload_0_2_2_6[7:0]   ), //i
    .push_payload_0_2_2_7     (streamDemux_2_io_outputs_7_payload_0_2_2_7[7:0]   ), //i
    .push_payload_0_2_2_8     (streamDemux_2_io_outputs_7_payload_0_2_2_8[7:0]   ), //i
    .push_payload_0_2_2_9     (streamDemux_2_io_outputs_7_payload_0_2_2_9[7:0]   ), //i
    .push_payload_0_2_2_10    (streamDemux_2_io_outputs_7_payload_0_2_2_10[7:0]  ), //i
    .push_payload_0_2_2_11    (streamDemux_2_io_outputs_7_payload_0_2_2_11[7:0]  ), //i
    .push_payload_0_2_2_12    (streamDemux_2_io_outputs_7_payload_0_2_2_12[7:0]  ), //i
    .push_payload_0_2_2_13    (streamDemux_2_io_outputs_7_payload_0_2_2_13[7:0]  ), //i
    .push_payload_0_2_2_14    (streamDemux_2_io_outputs_7_payload_0_2_2_14[7:0]  ), //i
    .push_payload_0_2_2_15    (streamDemux_2_io_outputs_7_payload_0_2_2_15[7:0]  ), //i
    .push_payload_1_0_0_0     (streamDemux_2_io_outputs_7_payload_1_0_0_0[7:0]   ), //i
    .push_payload_1_0_0_1     (streamDemux_2_io_outputs_7_payload_1_0_0_1[7:0]   ), //i
    .push_payload_1_0_0_2     (streamDemux_2_io_outputs_7_payload_1_0_0_2[7:0]   ), //i
    .push_payload_1_0_0_3     (streamDemux_2_io_outputs_7_payload_1_0_0_3[7:0]   ), //i
    .push_payload_1_0_0_4     (streamDemux_2_io_outputs_7_payload_1_0_0_4[7:0]   ), //i
    .push_payload_1_0_0_5     (streamDemux_2_io_outputs_7_payload_1_0_0_5[7:0]   ), //i
    .push_payload_1_0_0_6     (streamDemux_2_io_outputs_7_payload_1_0_0_6[7:0]   ), //i
    .push_payload_1_0_0_7     (streamDemux_2_io_outputs_7_payload_1_0_0_7[7:0]   ), //i
    .push_payload_1_0_0_8     (streamDemux_2_io_outputs_7_payload_1_0_0_8[7:0]   ), //i
    .push_payload_1_0_0_9     (streamDemux_2_io_outputs_7_payload_1_0_0_9[7:0]   ), //i
    .push_payload_1_0_0_10    (streamDemux_2_io_outputs_7_payload_1_0_0_10[7:0]  ), //i
    .push_payload_1_0_0_11    (streamDemux_2_io_outputs_7_payload_1_0_0_11[7:0]  ), //i
    .push_payload_1_0_0_12    (streamDemux_2_io_outputs_7_payload_1_0_0_12[7:0]  ), //i
    .push_payload_1_0_0_13    (streamDemux_2_io_outputs_7_payload_1_0_0_13[7:0]  ), //i
    .push_payload_1_0_0_14    (streamDemux_2_io_outputs_7_payload_1_0_0_14[7:0]  ), //i
    .push_payload_1_0_0_15    (streamDemux_2_io_outputs_7_payload_1_0_0_15[7:0]  ), //i
    .push_payload_1_0_1_0     (streamDemux_2_io_outputs_7_payload_1_0_1_0[7:0]   ), //i
    .push_payload_1_0_1_1     (streamDemux_2_io_outputs_7_payload_1_0_1_1[7:0]   ), //i
    .push_payload_1_0_1_2     (streamDemux_2_io_outputs_7_payload_1_0_1_2[7:0]   ), //i
    .push_payload_1_0_1_3     (streamDemux_2_io_outputs_7_payload_1_0_1_3[7:0]   ), //i
    .push_payload_1_0_1_4     (streamDemux_2_io_outputs_7_payload_1_0_1_4[7:0]   ), //i
    .push_payload_1_0_1_5     (streamDemux_2_io_outputs_7_payload_1_0_1_5[7:0]   ), //i
    .push_payload_1_0_1_6     (streamDemux_2_io_outputs_7_payload_1_0_1_6[7:0]   ), //i
    .push_payload_1_0_1_7     (streamDemux_2_io_outputs_7_payload_1_0_1_7[7:0]   ), //i
    .push_payload_1_0_1_8     (streamDemux_2_io_outputs_7_payload_1_0_1_8[7:0]   ), //i
    .push_payload_1_0_1_9     (streamDemux_2_io_outputs_7_payload_1_0_1_9[7:0]   ), //i
    .push_payload_1_0_1_10    (streamDemux_2_io_outputs_7_payload_1_0_1_10[7:0]  ), //i
    .push_payload_1_0_1_11    (streamDemux_2_io_outputs_7_payload_1_0_1_11[7:0]  ), //i
    .push_payload_1_0_1_12    (streamDemux_2_io_outputs_7_payload_1_0_1_12[7:0]  ), //i
    .push_payload_1_0_1_13    (streamDemux_2_io_outputs_7_payload_1_0_1_13[7:0]  ), //i
    .push_payload_1_0_1_14    (streamDemux_2_io_outputs_7_payload_1_0_1_14[7:0]  ), //i
    .push_payload_1_0_1_15    (streamDemux_2_io_outputs_7_payload_1_0_1_15[7:0]  ), //i
    .push_payload_1_0_2_0     (streamDemux_2_io_outputs_7_payload_1_0_2_0[7:0]   ), //i
    .push_payload_1_0_2_1     (streamDemux_2_io_outputs_7_payload_1_0_2_1[7:0]   ), //i
    .push_payload_1_0_2_2     (streamDemux_2_io_outputs_7_payload_1_0_2_2[7:0]   ), //i
    .push_payload_1_0_2_3     (streamDemux_2_io_outputs_7_payload_1_0_2_3[7:0]   ), //i
    .push_payload_1_0_2_4     (streamDemux_2_io_outputs_7_payload_1_0_2_4[7:0]   ), //i
    .push_payload_1_0_2_5     (streamDemux_2_io_outputs_7_payload_1_0_2_5[7:0]   ), //i
    .push_payload_1_0_2_6     (streamDemux_2_io_outputs_7_payload_1_0_2_6[7:0]   ), //i
    .push_payload_1_0_2_7     (streamDemux_2_io_outputs_7_payload_1_0_2_7[7:0]   ), //i
    .push_payload_1_0_2_8     (streamDemux_2_io_outputs_7_payload_1_0_2_8[7:0]   ), //i
    .push_payload_1_0_2_9     (streamDemux_2_io_outputs_7_payload_1_0_2_9[7:0]   ), //i
    .push_payload_1_0_2_10    (streamDemux_2_io_outputs_7_payload_1_0_2_10[7:0]  ), //i
    .push_payload_1_0_2_11    (streamDemux_2_io_outputs_7_payload_1_0_2_11[7:0]  ), //i
    .push_payload_1_0_2_12    (streamDemux_2_io_outputs_7_payload_1_0_2_12[7:0]  ), //i
    .push_payload_1_0_2_13    (streamDemux_2_io_outputs_7_payload_1_0_2_13[7:0]  ), //i
    .push_payload_1_0_2_14    (streamDemux_2_io_outputs_7_payload_1_0_2_14[7:0]  ), //i
    .push_payload_1_0_2_15    (streamDemux_2_io_outputs_7_payload_1_0_2_15[7:0]  ), //i
    .push_payload_1_1_0_0     (streamDemux_2_io_outputs_7_payload_1_1_0_0[7:0]   ), //i
    .push_payload_1_1_0_1     (streamDemux_2_io_outputs_7_payload_1_1_0_1[7:0]   ), //i
    .push_payload_1_1_0_2     (streamDemux_2_io_outputs_7_payload_1_1_0_2[7:0]   ), //i
    .push_payload_1_1_0_3     (streamDemux_2_io_outputs_7_payload_1_1_0_3[7:0]   ), //i
    .push_payload_1_1_0_4     (streamDemux_2_io_outputs_7_payload_1_1_0_4[7:0]   ), //i
    .push_payload_1_1_0_5     (streamDemux_2_io_outputs_7_payload_1_1_0_5[7:0]   ), //i
    .push_payload_1_1_0_6     (streamDemux_2_io_outputs_7_payload_1_1_0_6[7:0]   ), //i
    .push_payload_1_1_0_7     (streamDemux_2_io_outputs_7_payload_1_1_0_7[7:0]   ), //i
    .push_payload_1_1_0_8     (streamDemux_2_io_outputs_7_payload_1_1_0_8[7:0]   ), //i
    .push_payload_1_1_0_9     (streamDemux_2_io_outputs_7_payload_1_1_0_9[7:0]   ), //i
    .push_payload_1_1_0_10    (streamDemux_2_io_outputs_7_payload_1_1_0_10[7:0]  ), //i
    .push_payload_1_1_0_11    (streamDemux_2_io_outputs_7_payload_1_1_0_11[7:0]  ), //i
    .push_payload_1_1_0_12    (streamDemux_2_io_outputs_7_payload_1_1_0_12[7:0]  ), //i
    .push_payload_1_1_0_13    (streamDemux_2_io_outputs_7_payload_1_1_0_13[7:0]  ), //i
    .push_payload_1_1_0_14    (streamDemux_2_io_outputs_7_payload_1_1_0_14[7:0]  ), //i
    .push_payload_1_1_0_15    (streamDemux_2_io_outputs_7_payload_1_1_0_15[7:0]  ), //i
    .push_payload_1_1_1_0     (streamDemux_2_io_outputs_7_payload_1_1_1_0[7:0]   ), //i
    .push_payload_1_1_1_1     (streamDemux_2_io_outputs_7_payload_1_1_1_1[7:0]   ), //i
    .push_payload_1_1_1_2     (streamDemux_2_io_outputs_7_payload_1_1_1_2[7:0]   ), //i
    .push_payload_1_1_1_3     (streamDemux_2_io_outputs_7_payload_1_1_1_3[7:0]   ), //i
    .push_payload_1_1_1_4     (streamDemux_2_io_outputs_7_payload_1_1_1_4[7:0]   ), //i
    .push_payload_1_1_1_5     (streamDemux_2_io_outputs_7_payload_1_1_1_5[7:0]   ), //i
    .push_payload_1_1_1_6     (streamDemux_2_io_outputs_7_payload_1_1_1_6[7:0]   ), //i
    .push_payload_1_1_1_7     (streamDemux_2_io_outputs_7_payload_1_1_1_7[7:0]   ), //i
    .push_payload_1_1_1_8     (streamDemux_2_io_outputs_7_payload_1_1_1_8[7:0]   ), //i
    .push_payload_1_1_1_9     (streamDemux_2_io_outputs_7_payload_1_1_1_9[7:0]   ), //i
    .push_payload_1_1_1_10    (streamDemux_2_io_outputs_7_payload_1_1_1_10[7:0]  ), //i
    .push_payload_1_1_1_11    (streamDemux_2_io_outputs_7_payload_1_1_1_11[7:0]  ), //i
    .push_payload_1_1_1_12    (streamDemux_2_io_outputs_7_payload_1_1_1_12[7:0]  ), //i
    .push_payload_1_1_1_13    (streamDemux_2_io_outputs_7_payload_1_1_1_13[7:0]  ), //i
    .push_payload_1_1_1_14    (streamDemux_2_io_outputs_7_payload_1_1_1_14[7:0]  ), //i
    .push_payload_1_1_1_15    (streamDemux_2_io_outputs_7_payload_1_1_1_15[7:0]  ), //i
    .push_payload_1_1_2_0     (streamDemux_2_io_outputs_7_payload_1_1_2_0[7:0]   ), //i
    .push_payload_1_1_2_1     (streamDemux_2_io_outputs_7_payload_1_1_2_1[7:0]   ), //i
    .push_payload_1_1_2_2     (streamDemux_2_io_outputs_7_payload_1_1_2_2[7:0]   ), //i
    .push_payload_1_1_2_3     (streamDemux_2_io_outputs_7_payload_1_1_2_3[7:0]   ), //i
    .push_payload_1_1_2_4     (streamDemux_2_io_outputs_7_payload_1_1_2_4[7:0]   ), //i
    .push_payload_1_1_2_5     (streamDemux_2_io_outputs_7_payload_1_1_2_5[7:0]   ), //i
    .push_payload_1_1_2_6     (streamDemux_2_io_outputs_7_payload_1_1_2_6[7:0]   ), //i
    .push_payload_1_1_2_7     (streamDemux_2_io_outputs_7_payload_1_1_2_7[7:0]   ), //i
    .push_payload_1_1_2_8     (streamDemux_2_io_outputs_7_payload_1_1_2_8[7:0]   ), //i
    .push_payload_1_1_2_9     (streamDemux_2_io_outputs_7_payload_1_1_2_9[7:0]   ), //i
    .push_payload_1_1_2_10    (streamDemux_2_io_outputs_7_payload_1_1_2_10[7:0]  ), //i
    .push_payload_1_1_2_11    (streamDemux_2_io_outputs_7_payload_1_1_2_11[7:0]  ), //i
    .push_payload_1_1_2_12    (streamDemux_2_io_outputs_7_payload_1_1_2_12[7:0]  ), //i
    .push_payload_1_1_2_13    (streamDemux_2_io_outputs_7_payload_1_1_2_13[7:0]  ), //i
    .push_payload_1_1_2_14    (streamDemux_2_io_outputs_7_payload_1_1_2_14[7:0]  ), //i
    .push_payload_1_1_2_15    (streamDemux_2_io_outputs_7_payload_1_1_2_15[7:0]  ), //i
    .push_payload_1_2_0_0     (streamDemux_2_io_outputs_7_payload_1_2_0_0[7:0]   ), //i
    .push_payload_1_2_0_1     (streamDemux_2_io_outputs_7_payload_1_2_0_1[7:0]   ), //i
    .push_payload_1_2_0_2     (streamDemux_2_io_outputs_7_payload_1_2_0_2[7:0]   ), //i
    .push_payload_1_2_0_3     (streamDemux_2_io_outputs_7_payload_1_2_0_3[7:0]   ), //i
    .push_payload_1_2_0_4     (streamDemux_2_io_outputs_7_payload_1_2_0_4[7:0]   ), //i
    .push_payload_1_2_0_5     (streamDemux_2_io_outputs_7_payload_1_2_0_5[7:0]   ), //i
    .push_payload_1_2_0_6     (streamDemux_2_io_outputs_7_payload_1_2_0_6[7:0]   ), //i
    .push_payload_1_2_0_7     (streamDemux_2_io_outputs_7_payload_1_2_0_7[7:0]   ), //i
    .push_payload_1_2_0_8     (streamDemux_2_io_outputs_7_payload_1_2_0_8[7:0]   ), //i
    .push_payload_1_2_0_9     (streamDemux_2_io_outputs_7_payload_1_2_0_9[7:0]   ), //i
    .push_payload_1_2_0_10    (streamDemux_2_io_outputs_7_payload_1_2_0_10[7:0]  ), //i
    .push_payload_1_2_0_11    (streamDemux_2_io_outputs_7_payload_1_2_0_11[7:0]  ), //i
    .push_payload_1_2_0_12    (streamDemux_2_io_outputs_7_payload_1_2_0_12[7:0]  ), //i
    .push_payload_1_2_0_13    (streamDemux_2_io_outputs_7_payload_1_2_0_13[7:0]  ), //i
    .push_payload_1_2_0_14    (streamDemux_2_io_outputs_7_payload_1_2_0_14[7:0]  ), //i
    .push_payload_1_2_0_15    (streamDemux_2_io_outputs_7_payload_1_2_0_15[7:0]  ), //i
    .push_payload_1_2_1_0     (streamDemux_2_io_outputs_7_payload_1_2_1_0[7:0]   ), //i
    .push_payload_1_2_1_1     (streamDemux_2_io_outputs_7_payload_1_2_1_1[7:0]   ), //i
    .push_payload_1_2_1_2     (streamDemux_2_io_outputs_7_payload_1_2_1_2[7:0]   ), //i
    .push_payload_1_2_1_3     (streamDemux_2_io_outputs_7_payload_1_2_1_3[7:0]   ), //i
    .push_payload_1_2_1_4     (streamDemux_2_io_outputs_7_payload_1_2_1_4[7:0]   ), //i
    .push_payload_1_2_1_5     (streamDemux_2_io_outputs_7_payload_1_2_1_5[7:0]   ), //i
    .push_payload_1_2_1_6     (streamDemux_2_io_outputs_7_payload_1_2_1_6[7:0]   ), //i
    .push_payload_1_2_1_7     (streamDemux_2_io_outputs_7_payload_1_2_1_7[7:0]   ), //i
    .push_payload_1_2_1_8     (streamDemux_2_io_outputs_7_payload_1_2_1_8[7:0]   ), //i
    .push_payload_1_2_1_9     (streamDemux_2_io_outputs_7_payload_1_2_1_9[7:0]   ), //i
    .push_payload_1_2_1_10    (streamDemux_2_io_outputs_7_payload_1_2_1_10[7:0]  ), //i
    .push_payload_1_2_1_11    (streamDemux_2_io_outputs_7_payload_1_2_1_11[7:0]  ), //i
    .push_payload_1_2_1_12    (streamDemux_2_io_outputs_7_payload_1_2_1_12[7:0]  ), //i
    .push_payload_1_2_1_13    (streamDemux_2_io_outputs_7_payload_1_2_1_13[7:0]  ), //i
    .push_payload_1_2_1_14    (streamDemux_2_io_outputs_7_payload_1_2_1_14[7:0]  ), //i
    .push_payload_1_2_1_15    (streamDemux_2_io_outputs_7_payload_1_2_1_15[7:0]  ), //i
    .push_payload_1_2_2_0     (streamDemux_2_io_outputs_7_payload_1_2_2_0[7:0]   ), //i
    .push_payload_1_2_2_1     (streamDemux_2_io_outputs_7_payload_1_2_2_1[7:0]   ), //i
    .push_payload_1_2_2_2     (streamDemux_2_io_outputs_7_payload_1_2_2_2[7:0]   ), //i
    .push_payload_1_2_2_3     (streamDemux_2_io_outputs_7_payload_1_2_2_3[7:0]   ), //i
    .push_payload_1_2_2_4     (streamDemux_2_io_outputs_7_payload_1_2_2_4[7:0]   ), //i
    .push_payload_1_2_2_5     (streamDemux_2_io_outputs_7_payload_1_2_2_5[7:0]   ), //i
    .push_payload_1_2_2_6     (streamDemux_2_io_outputs_7_payload_1_2_2_6[7:0]   ), //i
    .push_payload_1_2_2_7     (streamDemux_2_io_outputs_7_payload_1_2_2_7[7:0]   ), //i
    .push_payload_1_2_2_8     (streamDemux_2_io_outputs_7_payload_1_2_2_8[7:0]   ), //i
    .push_payload_1_2_2_9     (streamDemux_2_io_outputs_7_payload_1_2_2_9[7:0]   ), //i
    .push_payload_1_2_2_10    (streamDemux_2_io_outputs_7_payload_1_2_2_10[7:0]  ), //i
    .push_payload_1_2_2_11    (streamDemux_2_io_outputs_7_payload_1_2_2_11[7:0]  ), //i
    .push_payload_1_2_2_12    (streamDemux_2_io_outputs_7_payload_1_2_2_12[7:0]  ), //i
    .push_payload_1_2_2_13    (streamDemux_2_io_outputs_7_payload_1_2_2_13[7:0]  ), //i
    .push_payload_1_2_2_14    (streamDemux_2_io_outputs_7_payload_1_2_2_14[7:0]  ), //i
    .push_payload_1_2_2_15    (streamDemux_2_io_outputs_7_payload_1_2_2_15[7:0]  ), //i
    .pop_valid                (weightFifo_7_pop_valid                            ), //o
    .pop_ready                (unit_7_weights_ready                              ), //i
    .pop_payload_0_0_0_0      (weightFifo_7_pop_payload_0_0_0_0[7:0]             ), //o
    .pop_payload_0_0_0_1      (weightFifo_7_pop_payload_0_0_0_1[7:0]             ), //o
    .pop_payload_0_0_0_2      (weightFifo_7_pop_payload_0_0_0_2[7:0]             ), //o
    .pop_payload_0_0_0_3      (weightFifo_7_pop_payload_0_0_0_3[7:0]             ), //o
    .pop_payload_0_0_0_4      (weightFifo_7_pop_payload_0_0_0_4[7:0]             ), //o
    .pop_payload_0_0_0_5      (weightFifo_7_pop_payload_0_0_0_5[7:0]             ), //o
    .pop_payload_0_0_0_6      (weightFifo_7_pop_payload_0_0_0_6[7:0]             ), //o
    .pop_payload_0_0_0_7      (weightFifo_7_pop_payload_0_0_0_7[7:0]             ), //o
    .pop_payload_0_0_0_8      (weightFifo_7_pop_payload_0_0_0_8[7:0]             ), //o
    .pop_payload_0_0_0_9      (weightFifo_7_pop_payload_0_0_0_9[7:0]             ), //o
    .pop_payload_0_0_0_10     (weightFifo_7_pop_payload_0_0_0_10[7:0]            ), //o
    .pop_payload_0_0_0_11     (weightFifo_7_pop_payload_0_0_0_11[7:0]            ), //o
    .pop_payload_0_0_0_12     (weightFifo_7_pop_payload_0_0_0_12[7:0]            ), //o
    .pop_payload_0_0_0_13     (weightFifo_7_pop_payload_0_0_0_13[7:0]            ), //o
    .pop_payload_0_0_0_14     (weightFifo_7_pop_payload_0_0_0_14[7:0]            ), //o
    .pop_payload_0_0_0_15     (weightFifo_7_pop_payload_0_0_0_15[7:0]            ), //o
    .pop_payload_0_0_1_0      (weightFifo_7_pop_payload_0_0_1_0[7:0]             ), //o
    .pop_payload_0_0_1_1      (weightFifo_7_pop_payload_0_0_1_1[7:0]             ), //o
    .pop_payload_0_0_1_2      (weightFifo_7_pop_payload_0_0_1_2[7:0]             ), //o
    .pop_payload_0_0_1_3      (weightFifo_7_pop_payload_0_0_1_3[7:0]             ), //o
    .pop_payload_0_0_1_4      (weightFifo_7_pop_payload_0_0_1_4[7:0]             ), //o
    .pop_payload_0_0_1_5      (weightFifo_7_pop_payload_0_0_1_5[7:0]             ), //o
    .pop_payload_0_0_1_6      (weightFifo_7_pop_payload_0_0_1_6[7:0]             ), //o
    .pop_payload_0_0_1_7      (weightFifo_7_pop_payload_0_0_1_7[7:0]             ), //o
    .pop_payload_0_0_1_8      (weightFifo_7_pop_payload_0_0_1_8[7:0]             ), //o
    .pop_payload_0_0_1_9      (weightFifo_7_pop_payload_0_0_1_9[7:0]             ), //o
    .pop_payload_0_0_1_10     (weightFifo_7_pop_payload_0_0_1_10[7:0]            ), //o
    .pop_payload_0_0_1_11     (weightFifo_7_pop_payload_0_0_1_11[7:0]            ), //o
    .pop_payload_0_0_1_12     (weightFifo_7_pop_payload_0_0_1_12[7:0]            ), //o
    .pop_payload_0_0_1_13     (weightFifo_7_pop_payload_0_0_1_13[7:0]            ), //o
    .pop_payload_0_0_1_14     (weightFifo_7_pop_payload_0_0_1_14[7:0]            ), //o
    .pop_payload_0_0_1_15     (weightFifo_7_pop_payload_0_0_1_15[7:0]            ), //o
    .pop_payload_0_0_2_0      (weightFifo_7_pop_payload_0_0_2_0[7:0]             ), //o
    .pop_payload_0_0_2_1      (weightFifo_7_pop_payload_0_0_2_1[7:0]             ), //o
    .pop_payload_0_0_2_2      (weightFifo_7_pop_payload_0_0_2_2[7:0]             ), //o
    .pop_payload_0_0_2_3      (weightFifo_7_pop_payload_0_0_2_3[7:0]             ), //o
    .pop_payload_0_0_2_4      (weightFifo_7_pop_payload_0_0_2_4[7:0]             ), //o
    .pop_payload_0_0_2_5      (weightFifo_7_pop_payload_0_0_2_5[7:0]             ), //o
    .pop_payload_0_0_2_6      (weightFifo_7_pop_payload_0_0_2_6[7:0]             ), //o
    .pop_payload_0_0_2_7      (weightFifo_7_pop_payload_0_0_2_7[7:0]             ), //o
    .pop_payload_0_0_2_8      (weightFifo_7_pop_payload_0_0_2_8[7:0]             ), //o
    .pop_payload_0_0_2_9      (weightFifo_7_pop_payload_0_0_2_9[7:0]             ), //o
    .pop_payload_0_0_2_10     (weightFifo_7_pop_payload_0_0_2_10[7:0]            ), //o
    .pop_payload_0_0_2_11     (weightFifo_7_pop_payload_0_0_2_11[7:0]            ), //o
    .pop_payload_0_0_2_12     (weightFifo_7_pop_payload_0_0_2_12[7:0]            ), //o
    .pop_payload_0_0_2_13     (weightFifo_7_pop_payload_0_0_2_13[7:0]            ), //o
    .pop_payload_0_0_2_14     (weightFifo_7_pop_payload_0_0_2_14[7:0]            ), //o
    .pop_payload_0_0_2_15     (weightFifo_7_pop_payload_0_0_2_15[7:0]            ), //o
    .pop_payload_0_1_0_0      (weightFifo_7_pop_payload_0_1_0_0[7:0]             ), //o
    .pop_payload_0_1_0_1      (weightFifo_7_pop_payload_0_1_0_1[7:0]             ), //o
    .pop_payload_0_1_0_2      (weightFifo_7_pop_payload_0_1_0_2[7:0]             ), //o
    .pop_payload_0_1_0_3      (weightFifo_7_pop_payload_0_1_0_3[7:0]             ), //o
    .pop_payload_0_1_0_4      (weightFifo_7_pop_payload_0_1_0_4[7:0]             ), //o
    .pop_payload_0_1_0_5      (weightFifo_7_pop_payload_0_1_0_5[7:0]             ), //o
    .pop_payload_0_1_0_6      (weightFifo_7_pop_payload_0_1_0_6[7:0]             ), //o
    .pop_payload_0_1_0_7      (weightFifo_7_pop_payload_0_1_0_7[7:0]             ), //o
    .pop_payload_0_1_0_8      (weightFifo_7_pop_payload_0_1_0_8[7:0]             ), //o
    .pop_payload_0_1_0_9      (weightFifo_7_pop_payload_0_1_0_9[7:0]             ), //o
    .pop_payload_0_1_0_10     (weightFifo_7_pop_payload_0_1_0_10[7:0]            ), //o
    .pop_payload_0_1_0_11     (weightFifo_7_pop_payload_0_1_0_11[7:0]            ), //o
    .pop_payload_0_1_0_12     (weightFifo_7_pop_payload_0_1_0_12[7:0]            ), //o
    .pop_payload_0_1_0_13     (weightFifo_7_pop_payload_0_1_0_13[7:0]            ), //o
    .pop_payload_0_1_0_14     (weightFifo_7_pop_payload_0_1_0_14[7:0]            ), //o
    .pop_payload_0_1_0_15     (weightFifo_7_pop_payload_0_1_0_15[7:0]            ), //o
    .pop_payload_0_1_1_0      (weightFifo_7_pop_payload_0_1_1_0[7:0]             ), //o
    .pop_payload_0_1_1_1      (weightFifo_7_pop_payload_0_1_1_1[7:0]             ), //o
    .pop_payload_0_1_1_2      (weightFifo_7_pop_payload_0_1_1_2[7:0]             ), //o
    .pop_payload_0_1_1_3      (weightFifo_7_pop_payload_0_1_1_3[7:0]             ), //o
    .pop_payload_0_1_1_4      (weightFifo_7_pop_payload_0_1_1_4[7:0]             ), //o
    .pop_payload_0_1_1_5      (weightFifo_7_pop_payload_0_1_1_5[7:0]             ), //o
    .pop_payload_0_1_1_6      (weightFifo_7_pop_payload_0_1_1_6[7:0]             ), //o
    .pop_payload_0_1_1_7      (weightFifo_7_pop_payload_0_1_1_7[7:0]             ), //o
    .pop_payload_0_1_1_8      (weightFifo_7_pop_payload_0_1_1_8[7:0]             ), //o
    .pop_payload_0_1_1_9      (weightFifo_7_pop_payload_0_1_1_9[7:0]             ), //o
    .pop_payload_0_1_1_10     (weightFifo_7_pop_payload_0_1_1_10[7:0]            ), //o
    .pop_payload_0_1_1_11     (weightFifo_7_pop_payload_0_1_1_11[7:0]            ), //o
    .pop_payload_0_1_1_12     (weightFifo_7_pop_payload_0_1_1_12[7:0]            ), //o
    .pop_payload_0_1_1_13     (weightFifo_7_pop_payload_0_1_1_13[7:0]            ), //o
    .pop_payload_0_1_1_14     (weightFifo_7_pop_payload_0_1_1_14[7:0]            ), //o
    .pop_payload_0_1_1_15     (weightFifo_7_pop_payload_0_1_1_15[7:0]            ), //o
    .pop_payload_0_1_2_0      (weightFifo_7_pop_payload_0_1_2_0[7:0]             ), //o
    .pop_payload_0_1_2_1      (weightFifo_7_pop_payload_0_1_2_1[7:0]             ), //o
    .pop_payload_0_1_2_2      (weightFifo_7_pop_payload_0_1_2_2[7:0]             ), //o
    .pop_payload_0_1_2_3      (weightFifo_7_pop_payload_0_1_2_3[7:0]             ), //o
    .pop_payload_0_1_2_4      (weightFifo_7_pop_payload_0_1_2_4[7:0]             ), //o
    .pop_payload_0_1_2_5      (weightFifo_7_pop_payload_0_1_2_5[7:0]             ), //o
    .pop_payload_0_1_2_6      (weightFifo_7_pop_payload_0_1_2_6[7:0]             ), //o
    .pop_payload_0_1_2_7      (weightFifo_7_pop_payload_0_1_2_7[7:0]             ), //o
    .pop_payload_0_1_2_8      (weightFifo_7_pop_payload_0_1_2_8[7:0]             ), //o
    .pop_payload_0_1_2_9      (weightFifo_7_pop_payload_0_1_2_9[7:0]             ), //o
    .pop_payload_0_1_2_10     (weightFifo_7_pop_payload_0_1_2_10[7:0]            ), //o
    .pop_payload_0_1_2_11     (weightFifo_7_pop_payload_0_1_2_11[7:0]            ), //o
    .pop_payload_0_1_2_12     (weightFifo_7_pop_payload_0_1_2_12[7:0]            ), //o
    .pop_payload_0_1_2_13     (weightFifo_7_pop_payload_0_1_2_13[7:0]            ), //o
    .pop_payload_0_1_2_14     (weightFifo_7_pop_payload_0_1_2_14[7:0]            ), //o
    .pop_payload_0_1_2_15     (weightFifo_7_pop_payload_0_1_2_15[7:0]            ), //o
    .pop_payload_0_2_0_0      (weightFifo_7_pop_payload_0_2_0_0[7:0]             ), //o
    .pop_payload_0_2_0_1      (weightFifo_7_pop_payload_0_2_0_1[7:0]             ), //o
    .pop_payload_0_2_0_2      (weightFifo_7_pop_payload_0_2_0_2[7:0]             ), //o
    .pop_payload_0_2_0_3      (weightFifo_7_pop_payload_0_2_0_3[7:0]             ), //o
    .pop_payload_0_2_0_4      (weightFifo_7_pop_payload_0_2_0_4[7:0]             ), //o
    .pop_payload_0_2_0_5      (weightFifo_7_pop_payload_0_2_0_5[7:0]             ), //o
    .pop_payload_0_2_0_6      (weightFifo_7_pop_payload_0_2_0_6[7:0]             ), //o
    .pop_payload_0_2_0_7      (weightFifo_7_pop_payload_0_2_0_7[7:0]             ), //o
    .pop_payload_0_2_0_8      (weightFifo_7_pop_payload_0_2_0_8[7:0]             ), //o
    .pop_payload_0_2_0_9      (weightFifo_7_pop_payload_0_2_0_9[7:0]             ), //o
    .pop_payload_0_2_0_10     (weightFifo_7_pop_payload_0_2_0_10[7:0]            ), //o
    .pop_payload_0_2_0_11     (weightFifo_7_pop_payload_0_2_0_11[7:0]            ), //o
    .pop_payload_0_2_0_12     (weightFifo_7_pop_payload_0_2_0_12[7:0]            ), //o
    .pop_payload_0_2_0_13     (weightFifo_7_pop_payload_0_2_0_13[7:0]            ), //o
    .pop_payload_0_2_0_14     (weightFifo_7_pop_payload_0_2_0_14[7:0]            ), //o
    .pop_payload_0_2_0_15     (weightFifo_7_pop_payload_0_2_0_15[7:0]            ), //o
    .pop_payload_0_2_1_0      (weightFifo_7_pop_payload_0_2_1_0[7:0]             ), //o
    .pop_payload_0_2_1_1      (weightFifo_7_pop_payload_0_2_1_1[7:0]             ), //o
    .pop_payload_0_2_1_2      (weightFifo_7_pop_payload_0_2_1_2[7:0]             ), //o
    .pop_payload_0_2_1_3      (weightFifo_7_pop_payload_0_2_1_3[7:0]             ), //o
    .pop_payload_0_2_1_4      (weightFifo_7_pop_payload_0_2_1_4[7:0]             ), //o
    .pop_payload_0_2_1_5      (weightFifo_7_pop_payload_0_2_1_5[7:0]             ), //o
    .pop_payload_0_2_1_6      (weightFifo_7_pop_payload_0_2_1_6[7:0]             ), //o
    .pop_payload_0_2_1_7      (weightFifo_7_pop_payload_0_2_1_7[7:0]             ), //o
    .pop_payload_0_2_1_8      (weightFifo_7_pop_payload_0_2_1_8[7:0]             ), //o
    .pop_payload_0_2_1_9      (weightFifo_7_pop_payload_0_2_1_9[7:0]             ), //o
    .pop_payload_0_2_1_10     (weightFifo_7_pop_payload_0_2_1_10[7:0]            ), //o
    .pop_payload_0_2_1_11     (weightFifo_7_pop_payload_0_2_1_11[7:0]            ), //o
    .pop_payload_0_2_1_12     (weightFifo_7_pop_payload_0_2_1_12[7:0]            ), //o
    .pop_payload_0_2_1_13     (weightFifo_7_pop_payload_0_2_1_13[7:0]            ), //o
    .pop_payload_0_2_1_14     (weightFifo_7_pop_payload_0_2_1_14[7:0]            ), //o
    .pop_payload_0_2_1_15     (weightFifo_7_pop_payload_0_2_1_15[7:0]            ), //o
    .pop_payload_0_2_2_0      (weightFifo_7_pop_payload_0_2_2_0[7:0]             ), //o
    .pop_payload_0_2_2_1      (weightFifo_7_pop_payload_0_2_2_1[7:0]             ), //o
    .pop_payload_0_2_2_2      (weightFifo_7_pop_payload_0_2_2_2[7:0]             ), //o
    .pop_payload_0_2_2_3      (weightFifo_7_pop_payload_0_2_2_3[7:0]             ), //o
    .pop_payload_0_2_2_4      (weightFifo_7_pop_payload_0_2_2_4[7:0]             ), //o
    .pop_payload_0_2_2_5      (weightFifo_7_pop_payload_0_2_2_5[7:0]             ), //o
    .pop_payload_0_2_2_6      (weightFifo_7_pop_payload_0_2_2_6[7:0]             ), //o
    .pop_payload_0_2_2_7      (weightFifo_7_pop_payload_0_2_2_7[7:0]             ), //o
    .pop_payload_0_2_2_8      (weightFifo_7_pop_payload_0_2_2_8[7:0]             ), //o
    .pop_payload_0_2_2_9      (weightFifo_7_pop_payload_0_2_2_9[7:0]             ), //o
    .pop_payload_0_2_2_10     (weightFifo_7_pop_payload_0_2_2_10[7:0]            ), //o
    .pop_payload_0_2_2_11     (weightFifo_7_pop_payload_0_2_2_11[7:0]            ), //o
    .pop_payload_0_2_2_12     (weightFifo_7_pop_payload_0_2_2_12[7:0]            ), //o
    .pop_payload_0_2_2_13     (weightFifo_7_pop_payload_0_2_2_13[7:0]            ), //o
    .pop_payload_0_2_2_14     (weightFifo_7_pop_payload_0_2_2_14[7:0]            ), //o
    .pop_payload_0_2_2_15     (weightFifo_7_pop_payload_0_2_2_15[7:0]            ), //o
    .pop_payload_1_0_0_0      (weightFifo_7_pop_payload_1_0_0_0[7:0]             ), //o
    .pop_payload_1_0_0_1      (weightFifo_7_pop_payload_1_0_0_1[7:0]             ), //o
    .pop_payload_1_0_0_2      (weightFifo_7_pop_payload_1_0_0_2[7:0]             ), //o
    .pop_payload_1_0_0_3      (weightFifo_7_pop_payload_1_0_0_3[7:0]             ), //o
    .pop_payload_1_0_0_4      (weightFifo_7_pop_payload_1_0_0_4[7:0]             ), //o
    .pop_payload_1_0_0_5      (weightFifo_7_pop_payload_1_0_0_5[7:0]             ), //o
    .pop_payload_1_0_0_6      (weightFifo_7_pop_payload_1_0_0_6[7:0]             ), //o
    .pop_payload_1_0_0_7      (weightFifo_7_pop_payload_1_0_0_7[7:0]             ), //o
    .pop_payload_1_0_0_8      (weightFifo_7_pop_payload_1_0_0_8[7:0]             ), //o
    .pop_payload_1_0_0_9      (weightFifo_7_pop_payload_1_0_0_9[7:0]             ), //o
    .pop_payload_1_0_0_10     (weightFifo_7_pop_payload_1_0_0_10[7:0]            ), //o
    .pop_payload_1_0_0_11     (weightFifo_7_pop_payload_1_0_0_11[7:0]            ), //o
    .pop_payload_1_0_0_12     (weightFifo_7_pop_payload_1_0_0_12[7:0]            ), //o
    .pop_payload_1_0_0_13     (weightFifo_7_pop_payload_1_0_0_13[7:0]            ), //o
    .pop_payload_1_0_0_14     (weightFifo_7_pop_payload_1_0_0_14[7:0]            ), //o
    .pop_payload_1_0_0_15     (weightFifo_7_pop_payload_1_0_0_15[7:0]            ), //o
    .pop_payload_1_0_1_0      (weightFifo_7_pop_payload_1_0_1_0[7:0]             ), //o
    .pop_payload_1_0_1_1      (weightFifo_7_pop_payload_1_0_1_1[7:0]             ), //o
    .pop_payload_1_0_1_2      (weightFifo_7_pop_payload_1_0_1_2[7:0]             ), //o
    .pop_payload_1_0_1_3      (weightFifo_7_pop_payload_1_0_1_3[7:0]             ), //o
    .pop_payload_1_0_1_4      (weightFifo_7_pop_payload_1_0_1_4[7:0]             ), //o
    .pop_payload_1_0_1_5      (weightFifo_7_pop_payload_1_0_1_5[7:0]             ), //o
    .pop_payload_1_0_1_6      (weightFifo_7_pop_payload_1_0_1_6[7:0]             ), //o
    .pop_payload_1_0_1_7      (weightFifo_7_pop_payload_1_0_1_7[7:0]             ), //o
    .pop_payload_1_0_1_8      (weightFifo_7_pop_payload_1_0_1_8[7:0]             ), //o
    .pop_payload_1_0_1_9      (weightFifo_7_pop_payload_1_0_1_9[7:0]             ), //o
    .pop_payload_1_0_1_10     (weightFifo_7_pop_payload_1_0_1_10[7:0]            ), //o
    .pop_payload_1_0_1_11     (weightFifo_7_pop_payload_1_0_1_11[7:0]            ), //o
    .pop_payload_1_0_1_12     (weightFifo_7_pop_payload_1_0_1_12[7:0]            ), //o
    .pop_payload_1_0_1_13     (weightFifo_7_pop_payload_1_0_1_13[7:0]            ), //o
    .pop_payload_1_0_1_14     (weightFifo_7_pop_payload_1_0_1_14[7:0]            ), //o
    .pop_payload_1_0_1_15     (weightFifo_7_pop_payload_1_0_1_15[7:0]            ), //o
    .pop_payload_1_0_2_0      (weightFifo_7_pop_payload_1_0_2_0[7:0]             ), //o
    .pop_payload_1_0_2_1      (weightFifo_7_pop_payload_1_0_2_1[7:0]             ), //o
    .pop_payload_1_0_2_2      (weightFifo_7_pop_payload_1_0_2_2[7:0]             ), //o
    .pop_payload_1_0_2_3      (weightFifo_7_pop_payload_1_0_2_3[7:0]             ), //o
    .pop_payload_1_0_2_4      (weightFifo_7_pop_payload_1_0_2_4[7:0]             ), //o
    .pop_payload_1_0_2_5      (weightFifo_7_pop_payload_1_0_2_5[7:0]             ), //o
    .pop_payload_1_0_2_6      (weightFifo_7_pop_payload_1_0_2_6[7:0]             ), //o
    .pop_payload_1_0_2_7      (weightFifo_7_pop_payload_1_0_2_7[7:0]             ), //o
    .pop_payload_1_0_2_8      (weightFifo_7_pop_payload_1_0_2_8[7:0]             ), //o
    .pop_payload_1_0_2_9      (weightFifo_7_pop_payload_1_0_2_9[7:0]             ), //o
    .pop_payload_1_0_2_10     (weightFifo_7_pop_payload_1_0_2_10[7:0]            ), //o
    .pop_payload_1_0_2_11     (weightFifo_7_pop_payload_1_0_2_11[7:0]            ), //o
    .pop_payload_1_0_2_12     (weightFifo_7_pop_payload_1_0_2_12[7:0]            ), //o
    .pop_payload_1_0_2_13     (weightFifo_7_pop_payload_1_0_2_13[7:0]            ), //o
    .pop_payload_1_0_2_14     (weightFifo_7_pop_payload_1_0_2_14[7:0]            ), //o
    .pop_payload_1_0_2_15     (weightFifo_7_pop_payload_1_0_2_15[7:0]            ), //o
    .pop_payload_1_1_0_0      (weightFifo_7_pop_payload_1_1_0_0[7:0]             ), //o
    .pop_payload_1_1_0_1      (weightFifo_7_pop_payload_1_1_0_1[7:0]             ), //o
    .pop_payload_1_1_0_2      (weightFifo_7_pop_payload_1_1_0_2[7:0]             ), //o
    .pop_payload_1_1_0_3      (weightFifo_7_pop_payload_1_1_0_3[7:0]             ), //o
    .pop_payload_1_1_0_4      (weightFifo_7_pop_payload_1_1_0_4[7:0]             ), //o
    .pop_payload_1_1_0_5      (weightFifo_7_pop_payload_1_1_0_5[7:0]             ), //o
    .pop_payload_1_1_0_6      (weightFifo_7_pop_payload_1_1_0_6[7:0]             ), //o
    .pop_payload_1_1_0_7      (weightFifo_7_pop_payload_1_1_0_7[7:0]             ), //o
    .pop_payload_1_1_0_8      (weightFifo_7_pop_payload_1_1_0_8[7:0]             ), //o
    .pop_payload_1_1_0_9      (weightFifo_7_pop_payload_1_1_0_9[7:0]             ), //o
    .pop_payload_1_1_0_10     (weightFifo_7_pop_payload_1_1_0_10[7:0]            ), //o
    .pop_payload_1_1_0_11     (weightFifo_7_pop_payload_1_1_0_11[7:0]            ), //o
    .pop_payload_1_1_0_12     (weightFifo_7_pop_payload_1_1_0_12[7:0]            ), //o
    .pop_payload_1_1_0_13     (weightFifo_7_pop_payload_1_1_0_13[7:0]            ), //o
    .pop_payload_1_1_0_14     (weightFifo_7_pop_payload_1_1_0_14[7:0]            ), //o
    .pop_payload_1_1_0_15     (weightFifo_7_pop_payload_1_1_0_15[7:0]            ), //o
    .pop_payload_1_1_1_0      (weightFifo_7_pop_payload_1_1_1_0[7:0]             ), //o
    .pop_payload_1_1_1_1      (weightFifo_7_pop_payload_1_1_1_1[7:0]             ), //o
    .pop_payload_1_1_1_2      (weightFifo_7_pop_payload_1_1_1_2[7:0]             ), //o
    .pop_payload_1_1_1_3      (weightFifo_7_pop_payload_1_1_1_3[7:0]             ), //o
    .pop_payload_1_1_1_4      (weightFifo_7_pop_payload_1_1_1_4[7:0]             ), //o
    .pop_payload_1_1_1_5      (weightFifo_7_pop_payload_1_1_1_5[7:0]             ), //o
    .pop_payload_1_1_1_6      (weightFifo_7_pop_payload_1_1_1_6[7:0]             ), //o
    .pop_payload_1_1_1_7      (weightFifo_7_pop_payload_1_1_1_7[7:0]             ), //o
    .pop_payload_1_1_1_8      (weightFifo_7_pop_payload_1_1_1_8[7:0]             ), //o
    .pop_payload_1_1_1_9      (weightFifo_7_pop_payload_1_1_1_9[7:0]             ), //o
    .pop_payload_1_1_1_10     (weightFifo_7_pop_payload_1_1_1_10[7:0]            ), //o
    .pop_payload_1_1_1_11     (weightFifo_7_pop_payload_1_1_1_11[7:0]            ), //o
    .pop_payload_1_1_1_12     (weightFifo_7_pop_payload_1_1_1_12[7:0]            ), //o
    .pop_payload_1_1_1_13     (weightFifo_7_pop_payload_1_1_1_13[7:0]            ), //o
    .pop_payload_1_1_1_14     (weightFifo_7_pop_payload_1_1_1_14[7:0]            ), //o
    .pop_payload_1_1_1_15     (weightFifo_7_pop_payload_1_1_1_15[7:0]            ), //o
    .pop_payload_1_1_2_0      (weightFifo_7_pop_payload_1_1_2_0[7:0]             ), //o
    .pop_payload_1_1_2_1      (weightFifo_7_pop_payload_1_1_2_1[7:0]             ), //o
    .pop_payload_1_1_2_2      (weightFifo_7_pop_payload_1_1_2_2[7:0]             ), //o
    .pop_payload_1_1_2_3      (weightFifo_7_pop_payload_1_1_2_3[7:0]             ), //o
    .pop_payload_1_1_2_4      (weightFifo_7_pop_payload_1_1_2_4[7:0]             ), //o
    .pop_payload_1_1_2_5      (weightFifo_7_pop_payload_1_1_2_5[7:0]             ), //o
    .pop_payload_1_1_2_6      (weightFifo_7_pop_payload_1_1_2_6[7:0]             ), //o
    .pop_payload_1_1_2_7      (weightFifo_7_pop_payload_1_1_2_7[7:0]             ), //o
    .pop_payload_1_1_2_8      (weightFifo_7_pop_payload_1_1_2_8[7:0]             ), //o
    .pop_payload_1_1_2_9      (weightFifo_7_pop_payload_1_1_2_9[7:0]             ), //o
    .pop_payload_1_1_2_10     (weightFifo_7_pop_payload_1_1_2_10[7:0]            ), //o
    .pop_payload_1_1_2_11     (weightFifo_7_pop_payload_1_1_2_11[7:0]            ), //o
    .pop_payload_1_1_2_12     (weightFifo_7_pop_payload_1_1_2_12[7:0]            ), //o
    .pop_payload_1_1_2_13     (weightFifo_7_pop_payload_1_1_2_13[7:0]            ), //o
    .pop_payload_1_1_2_14     (weightFifo_7_pop_payload_1_1_2_14[7:0]            ), //o
    .pop_payload_1_1_2_15     (weightFifo_7_pop_payload_1_1_2_15[7:0]            ), //o
    .pop_payload_1_2_0_0      (weightFifo_7_pop_payload_1_2_0_0[7:0]             ), //o
    .pop_payload_1_2_0_1      (weightFifo_7_pop_payload_1_2_0_1[7:0]             ), //o
    .pop_payload_1_2_0_2      (weightFifo_7_pop_payload_1_2_0_2[7:0]             ), //o
    .pop_payload_1_2_0_3      (weightFifo_7_pop_payload_1_2_0_3[7:0]             ), //o
    .pop_payload_1_2_0_4      (weightFifo_7_pop_payload_1_2_0_4[7:0]             ), //o
    .pop_payload_1_2_0_5      (weightFifo_7_pop_payload_1_2_0_5[7:0]             ), //o
    .pop_payload_1_2_0_6      (weightFifo_7_pop_payload_1_2_0_6[7:0]             ), //o
    .pop_payload_1_2_0_7      (weightFifo_7_pop_payload_1_2_0_7[7:0]             ), //o
    .pop_payload_1_2_0_8      (weightFifo_7_pop_payload_1_2_0_8[7:0]             ), //o
    .pop_payload_1_2_0_9      (weightFifo_7_pop_payload_1_2_0_9[7:0]             ), //o
    .pop_payload_1_2_0_10     (weightFifo_7_pop_payload_1_2_0_10[7:0]            ), //o
    .pop_payload_1_2_0_11     (weightFifo_7_pop_payload_1_2_0_11[7:0]            ), //o
    .pop_payload_1_2_0_12     (weightFifo_7_pop_payload_1_2_0_12[7:0]            ), //o
    .pop_payload_1_2_0_13     (weightFifo_7_pop_payload_1_2_0_13[7:0]            ), //o
    .pop_payload_1_2_0_14     (weightFifo_7_pop_payload_1_2_0_14[7:0]            ), //o
    .pop_payload_1_2_0_15     (weightFifo_7_pop_payload_1_2_0_15[7:0]            ), //o
    .pop_payload_1_2_1_0      (weightFifo_7_pop_payload_1_2_1_0[7:0]             ), //o
    .pop_payload_1_2_1_1      (weightFifo_7_pop_payload_1_2_1_1[7:0]             ), //o
    .pop_payload_1_2_1_2      (weightFifo_7_pop_payload_1_2_1_2[7:0]             ), //o
    .pop_payload_1_2_1_3      (weightFifo_7_pop_payload_1_2_1_3[7:0]             ), //o
    .pop_payload_1_2_1_4      (weightFifo_7_pop_payload_1_2_1_4[7:0]             ), //o
    .pop_payload_1_2_1_5      (weightFifo_7_pop_payload_1_2_1_5[7:0]             ), //o
    .pop_payload_1_2_1_6      (weightFifo_7_pop_payload_1_2_1_6[7:0]             ), //o
    .pop_payload_1_2_1_7      (weightFifo_7_pop_payload_1_2_1_7[7:0]             ), //o
    .pop_payload_1_2_1_8      (weightFifo_7_pop_payload_1_2_1_8[7:0]             ), //o
    .pop_payload_1_2_1_9      (weightFifo_7_pop_payload_1_2_1_9[7:0]             ), //o
    .pop_payload_1_2_1_10     (weightFifo_7_pop_payload_1_2_1_10[7:0]            ), //o
    .pop_payload_1_2_1_11     (weightFifo_7_pop_payload_1_2_1_11[7:0]            ), //o
    .pop_payload_1_2_1_12     (weightFifo_7_pop_payload_1_2_1_12[7:0]            ), //o
    .pop_payload_1_2_1_13     (weightFifo_7_pop_payload_1_2_1_13[7:0]            ), //o
    .pop_payload_1_2_1_14     (weightFifo_7_pop_payload_1_2_1_14[7:0]            ), //o
    .pop_payload_1_2_1_15     (weightFifo_7_pop_payload_1_2_1_15[7:0]            ), //o
    .pop_payload_1_2_2_0      (weightFifo_7_pop_payload_1_2_2_0[7:0]             ), //o
    .pop_payload_1_2_2_1      (weightFifo_7_pop_payload_1_2_2_1[7:0]             ), //o
    .pop_payload_1_2_2_2      (weightFifo_7_pop_payload_1_2_2_2[7:0]             ), //o
    .pop_payload_1_2_2_3      (weightFifo_7_pop_payload_1_2_2_3[7:0]             ), //o
    .pop_payload_1_2_2_4      (weightFifo_7_pop_payload_1_2_2_4[7:0]             ), //o
    .pop_payload_1_2_2_5      (weightFifo_7_pop_payload_1_2_2_5[7:0]             ), //o
    .pop_payload_1_2_2_6      (weightFifo_7_pop_payload_1_2_2_6[7:0]             ), //o
    .pop_payload_1_2_2_7      (weightFifo_7_pop_payload_1_2_2_7[7:0]             ), //o
    .pop_payload_1_2_2_8      (weightFifo_7_pop_payload_1_2_2_8[7:0]             ), //o
    .pop_payload_1_2_2_9      (weightFifo_7_pop_payload_1_2_2_9[7:0]             ), //o
    .pop_payload_1_2_2_10     (weightFifo_7_pop_payload_1_2_2_10[7:0]            ), //o
    .pop_payload_1_2_2_11     (weightFifo_7_pop_payload_1_2_2_11[7:0]            ), //o
    .pop_payload_1_2_2_12     (weightFifo_7_pop_payload_1_2_2_12[7:0]            ), //o
    .pop_payload_1_2_2_13     (weightFifo_7_pop_payload_1_2_2_13[7:0]            ), //o
    .pop_payload_1_2_2_14     (weightFifo_7_pop_payload_1_2_2_14[7:0]            ), //o
    .pop_payload_1_2_2_15     (weightFifo_7_pop_payload_1_2_2_15[7:0]            ), //o
    .flush                    (1'b0                                              ), //i
    .clk                      (clk                                               ), //i
    .reset                    (reset                                             )  //i
  );
  SlidingWindowSame window (
    .videoIn_valid                               (inputVideo_valid                                      ), //i
    .videoIn_ready                               (window_videoIn_ready                                  ), //o
    .videoIn_payload_frame_line_pixel_0          (inputVideo_payload_frame_line_pixel_0[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_1          (inputVideo_payload_frame_line_pixel_1[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_2          (inputVideo_payload_frame_line_pixel_2[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_3          (inputVideo_payload_frame_line_pixel_3[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_4          (inputVideo_payload_frame_line_pixel_4[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_5          (inputVideo_payload_frame_line_pixel_5[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_6          (inputVideo_payload_frame_line_pixel_6[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_7          (inputVideo_payload_frame_line_pixel_7[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_8          (inputVideo_payload_frame_line_pixel_8[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_9          (inputVideo_payload_frame_line_pixel_9[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_10         (inputVideo_payload_frame_line_pixel_10[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_11         (inputVideo_payload_frame_line_pixel_11[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_12         (inputVideo_payload_frame_line_pixel_12[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_13         (inputVideo_payload_frame_line_pixel_13[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_14         (inputVideo_payload_frame_line_pixel_14[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_15         (inputVideo_payload_frame_line_pixel_15[7:0]           ), //i
    .videoIn_payload_frame_line_endOfLine        (inputVideo_payload_frame_line_endOfLine               ), //i
    .videoIn_payload_frame_endOfFrame            (inputVideo_payload_frame_endOfFrame                   ), //i
    .videoIn_payload_endOfPack                   (inputVideo_payload_endOfPack                          ), //i
    .videoOut_valid                              (window_videoOut_valid                                 ), //o
    .videoOut_ready                              (window_videoOut_fork_io_input_ready                   ), //i
    .videoOut_payload_frame_line_pixel_0_0_0     (window_videoOut_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_1     (window_videoOut_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_2     (window_videoOut_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_3     (window_videoOut_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_4     (window_videoOut_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_5     (window_videoOut_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_6     (window_videoOut_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_7     (window_videoOut_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_8     (window_videoOut_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_9     (window_videoOut_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_10    (window_videoOut_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_11    (window_videoOut_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_12    (window_videoOut_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_13    (window_videoOut_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_14    (window_videoOut_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_15    (window_videoOut_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_0     (window_videoOut_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_1     (window_videoOut_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_2     (window_videoOut_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_3     (window_videoOut_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_4     (window_videoOut_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_5     (window_videoOut_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_6     (window_videoOut_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_7     (window_videoOut_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_8     (window_videoOut_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_9     (window_videoOut_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_10    (window_videoOut_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_11    (window_videoOut_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_12    (window_videoOut_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_13    (window_videoOut_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_14    (window_videoOut_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_15    (window_videoOut_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_0     (window_videoOut_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_1     (window_videoOut_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_2     (window_videoOut_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_3     (window_videoOut_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_4     (window_videoOut_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_5     (window_videoOut_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_6     (window_videoOut_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_7     (window_videoOut_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_8     (window_videoOut_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_9     (window_videoOut_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2_10    (window_videoOut_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_11    (window_videoOut_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_12    (window_videoOut_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_13    (window_videoOut_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_14    (window_videoOut_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_2_15    (window_videoOut_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_0     (window_videoOut_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_1     (window_videoOut_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_2     (window_videoOut_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_3     (window_videoOut_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_4     (window_videoOut_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_5     (window_videoOut_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_6     (window_videoOut_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_7     (window_videoOut_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_8     (window_videoOut_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_9     (window_videoOut_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_10    (window_videoOut_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_11    (window_videoOut_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_12    (window_videoOut_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_13    (window_videoOut_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_14    (window_videoOut_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_15    (window_videoOut_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_0     (window_videoOut_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_1     (window_videoOut_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_2     (window_videoOut_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_3     (window_videoOut_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_4     (window_videoOut_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_5     (window_videoOut_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_6     (window_videoOut_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_7     (window_videoOut_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_8     (window_videoOut_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_9     (window_videoOut_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_10    (window_videoOut_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_11    (window_videoOut_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_12    (window_videoOut_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_13    (window_videoOut_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_14    (window_videoOut_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_15    (window_videoOut_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_0     (window_videoOut_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_1     (window_videoOut_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_2     (window_videoOut_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_3     (window_videoOut_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_4     (window_videoOut_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_5     (window_videoOut_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_6     (window_videoOut_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_7     (window_videoOut_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_8     (window_videoOut_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_9     (window_videoOut_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2_10    (window_videoOut_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_11    (window_videoOut_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_12    (window_videoOut_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_13    (window_videoOut_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_14    (window_videoOut_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_2_15    (window_videoOut_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_0     (window_videoOut_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_1     (window_videoOut_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_2     (window_videoOut_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_3     (window_videoOut_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_4     (window_videoOut_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_5     (window_videoOut_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_6     (window_videoOut_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_7     (window_videoOut_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_8     (window_videoOut_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_9     (window_videoOut_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_0_10    (window_videoOut_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_11    (window_videoOut_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_12    (window_videoOut_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_13    (window_videoOut_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_14    (window_videoOut_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0_15    (window_videoOut_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_0     (window_videoOut_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_1     (window_videoOut_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_2     (window_videoOut_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_3     (window_videoOut_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_4     (window_videoOut_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_5     (window_videoOut_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_6     (window_videoOut_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_7     (window_videoOut_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_8     (window_videoOut_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_9     (window_videoOut_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1_10    (window_videoOut_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_11    (window_videoOut_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_12    (window_videoOut_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_13    (window_videoOut_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_14    (window_videoOut_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_1_15    (window_videoOut_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_0     (window_videoOut_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_1     (window_videoOut_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_2     (window_videoOut_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_3     (window_videoOut_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_4     (window_videoOut_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_5     (window_videoOut_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_6     (window_videoOut_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_7     (window_videoOut_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_8     (window_videoOut_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_9     (window_videoOut_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2_10    (window_videoOut_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_11    (window_videoOut_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_12    (window_videoOut_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_13    (window_videoOut_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_14    (window_videoOut_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_2_15    (window_videoOut_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .videoOut_payload_frame_line_endOfLine       (window_videoOut_payload_frame_line_endOfLine          ), //o
    .videoOut_payload_frame_endOfFrame           (window_videoOut_payload_frame_endOfFrame              ), //o
    .videoOut_payload_endOfPack                  (window_videoOut_payload_endOfPack                     ), //o
    .clk                                         (clk                                                   ), //i
    .reset                                       (reset                                                 )  //i
  );
  StreamFork_4 window_videoOut_fork (
    .io_input_valid                                  (window_videoOut_valid                                                   ), //i
    .io_input_ready                                  (window_videoOut_fork_io_input_ready                                     ), //o
    .io_input_payload_frame_line_pixel_0_0_0         (window_videoOut_payload_frame_line_pixel_0_0_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_1         (window_videoOut_payload_frame_line_pixel_0_0_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_2         (window_videoOut_payload_frame_line_pixel_0_0_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_3         (window_videoOut_payload_frame_line_pixel_0_0_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_4         (window_videoOut_payload_frame_line_pixel_0_0_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_5         (window_videoOut_payload_frame_line_pixel_0_0_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_6         (window_videoOut_payload_frame_line_pixel_0_0_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_7         (window_videoOut_payload_frame_line_pixel_0_0_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_8         (window_videoOut_payload_frame_line_pixel_0_0_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_9         (window_videoOut_payload_frame_line_pixel_0_0_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_0_10        (window_videoOut_payload_frame_line_pixel_0_0_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_0_11        (window_videoOut_payload_frame_line_pixel_0_0_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_0_12        (window_videoOut_payload_frame_line_pixel_0_0_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_0_13        (window_videoOut_payload_frame_line_pixel_0_0_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_0_14        (window_videoOut_payload_frame_line_pixel_0_0_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_0_15        (window_videoOut_payload_frame_line_pixel_0_0_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_0         (window_videoOut_payload_frame_line_pixel_0_1_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_1         (window_videoOut_payload_frame_line_pixel_0_1_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_2         (window_videoOut_payload_frame_line_pixel_0_1_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_3         (window_videoOut_payload_frame_line_pixel_0_1_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_4         (window_videoOut_payload_frame_line_pixel_0_1_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_5         (window_videoOut_payload_frame_line_pixel_0_1_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_6         (window_videoOut_payload_frame_line_pixel_0_1_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_7         (window_videoOut_payload_frame_line_pixel_0_1_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_8         (window_videoOut_payload_frame_line_pixel_0_1_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_9         (window_videoOut_payload_frame_line_pixel_0_1_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_1_10        (window_videoOut_payload_frame_line_pixel_0_1_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_11        (window_videoOut_payload_frame_line_pixel_0_1_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_12        (window_videoOut_payload_frame_line_pixel_0_1_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_13        (window_videoOut_payload_frame_line_pixel_0_1_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_14        (window_videoOut_payload_frame_line_pixel_0_1_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_1_15        (window_videoOut_payload_frame_line_pixel_0_1_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_0         (window_videoOut_payload_frame_line_pixel_0_2_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_1         (window_videoOut_payload_frame_line_pixel_0_2_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_2         (window_videoOut_payload_frame_line_pixel_0_2_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_3         (window_videoOut_payload_frame_line_pixel_0_2_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_4         (window_videoOut_payload_frame_line_pixel_0_2_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_5         (window_videoOut_payload_frame_line_pixel_0_2_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_6         (window_videoOut_payload_frame_line_pixel_0_2_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_7         (window_videoOut_payload_frame_line_pixel_0_2_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_8         (window_videoOut_payload_frame_line_pixel_0_2_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_9         (window_videoOut_payload_frame_line_pixel_0_2_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_0_2_10        (window_videoOut_payload_frame_line_pixel_0_2_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_11        (window_videoOut_payload_frame_line_pixel_0_2_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_12        (window_videoOut_payload_frame_line_pixel_0_2_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_13        (window_videoOut_payload_frame_line_pixel_0_2_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_14        (window_videoOut_payload_frame_line_pixel_0_2_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_0_2_15        (window_videoOut_payload_frame_line_pixel_0_2_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_0         (window_videoOut_payload_frame_line_pixel_1_0_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_1         (window_videoOut_payload_frame_line_pixel_1_0_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_2         (window_videoOut_payload_frame_line_pixel_1_0_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_3         (window_videoOut_payload_frame_line_pixel_1_0_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_4         (window_videoOut_payload_frame_line_pixel_1_0_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_5         (window_videoOut_payload_frame_line_pixel_1_0_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_6         (window_videoOut_payload_frame_line_pixel_1_0_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_7         (window_videoOut_payload_frame_line_pixel_1_0_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_8         (window_videoOut_payload_frame_line_pixel_1_0_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_9         (window_videoOut_payload_frame_line_pixel_1_0_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_0_10        (window_videoOut_payload_frame_line_pixel_1_0_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_11        (window_videoOut_payload_frame_line_pixel_1_0_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_12        (window_videoOut_payload_frame_line_pixel_1_0_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_13        (window_videoOut_payload_frame_line_pixel_1_0_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_14        (window_videoOut_payload_frame_line_pixel_1_0_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_0_15        (window_videoOut_payload_frame_line_pixel_1_0_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_0         (window_videoOut_payload_frame_line_pixel_1_1_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_1         (window_videoOut_payload_frame_line_pixel_1_1_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_2         (window_videoOut_payload_frame_line_pixel_1_1_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_3         (window_videoOut_payload_frame_line_pixel_1_1_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_4         (window_videoOut_payload_frame_line_pixel_1_1_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_5         (window_videoOut_payload_frame_line_pixel_1_1_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_6         (window_videoOut_payload_frame_line_pixel_1_1_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_7         (window_videoOut_payload_frame_line_pixel_1_1_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_8         (window_videoOut_payload_frame_line_pixel_1_1_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_9         (window_videoOut_payload_frame_line_pixel_1_1_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_1_10        (window_videoOut_payload_frame_line_pixel_1_1_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_11        (window_videoOut_payload_frame_line_pixel_1_1_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_12        (window_videoOut_payload_frame_line_pixel_1_1_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_13        (window_videoOut_payload_frame_line_pixel_1_1_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_14        (window_videoOut_payload_frame_line_pixel_1_1_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_1_15        (window_videoOut_payload_frame_line_pixel_1_1_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_0         (window_videoOut_payload_frame_line_pixel_1_2_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_1         (window_videoOut_payload_frame_line_pixel_1_2_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_2         (window_videoOut_payload_frame_line_pixel_1_2_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_3         (window_videoOut_payload_frame_line_pixel_1_2_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_4         (window_videoOut_payload_frame_line_pixel_1_2_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_5         (window_videoOut_payload_frame_line_pixel_1_2_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_6         (window_videoOut_payload_frame_line_pixel_1_2_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_7         (window_videoOut_payload_frame_line_pixel_1_2_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_8         (window_videoOut_payload_frame_line_pixel_1_2_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_9         (window_videoOut_payload_frame_line_pixel_1_2_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1_2_10        (window_videoOut_payload_frame_line_pixel_1_2_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_11        (window_videoOut_payload_frame_line_pixel_1_2_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_12        (window_videoOut_payload_frame_line_pixel_1_2_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_13        (window_videoOut_payload_frame_line_pixel_1_2_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_14        (window_videoOut_payload_frame_line_pixel_1_2_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_1_2_15        (window_videoOut_payload_frame_line_pixel_1_2_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_0         (window_videoOut_payload_frame_line_pixel_2_0_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_1         (window_videoOut_payload_frame_line_pixel_2_0_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_2         (window_videoOut_payload_frame_line_pixel_2_0_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_3         (window_videoOut_payload_frame_line_pixel_2_0_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_4         (window_videoOut_payload_frame_line_pixel_2_0_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_5         (window_videoOut_payload_frame_line_pixel_2_0_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_6         (window_videoOut_payload_frame_line_pixel_2_0_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_7         (window_videoOut_payload_frame_line_pixel_2_0_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_8         (window_videoOut_payload_frame_line_pixel_2_0_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_9         (window_videoOut_payload_frame_line_pixel_2_0_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_0_10        (window_videoOut_payload_frame_line_pixel_2_0_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_11        (window_videoOut_payload_frame_line_pixel_2_0_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_12        (window_videoOut_payload_frame_line_pixel_2_0_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_13        (window_videoOut_payload_frame_line_pixel_2_0_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_14        (window_videoOut_payload_frame_line_pixel_2_0_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_0_15        (window_videoOut_payload_frame_line_pixel_2_0_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_0         (window_videoOut_payload_frame_line_pixel_2_1_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_1         (window_videoOut_payload_frame_line_pixel_2_1_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_2         (window_videoOut_payload_frame_line_pixel_2_1_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_3         (window_videoOut_payload_frame_line_pixel_2_1_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_4         (window_videoOut_payload_frame_line_pixel_2_1_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_5         (window_videoOut_payload_frame_line_pixel_2_1_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_6         (window_videoOut_payload_frame_line_pixel_2_1_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_7         (window_videoOut_payload_frame_line_pixel_2_1_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_8         (window_videoOut_payload_frame_line_pixel_2_1_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_9         (window_videoOut_payload_frame_line_pixel_2_1_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_1_10        (window_videoOut_payload_frame_line_pixel_2_1_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_11        (window_videoOut_payload_frame_line_pixel_2_1_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_12        (window_videoOut_payload_frame_line_pixel_2_1_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_13        (window_videoOut_payload_frame_line_pixel_2_1_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_14        (window_videoOut_payload_frame_line_pixel_2_1_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_1_15        (window_videoOut_payload_frame_line_pixel_2_1_15[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_0         (window_videoOut_payload_frame_line_pixel_2_2_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_1         (window_videoOut_payload_frame_line_pixel_2_2_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_2         (window_videoOut_payload_frame_line_pixel_2_2_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_3         (window_videoOut_payload_frame_line_pixel_2_2_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_4         (window_videoOut_payload_frame_line_pixel_2_2_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_5         (window_videoOut_payload_frame_line_pixel_2_2_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_6         (window_videoOut_payload_frame_line_pixel_2_2_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_7         (window_videoOut_payload_frame_line_pixel_2_2_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_8         (window_videoOut_payload_frame_line_pixel_2_2_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_9         (window_videoOut_payload_frame_line_pixel_2_2_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2_2_10        (window_videoOut_payload_frame_line_pixel_2_2_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_11        (window_videoOut_payload_frame_line_pixel_2_2_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_12        (window_videoOut_payload_frame_line_pixel_2_2_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_13        (window_videoOut_payload_frame_line_pixel_2_2_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_14        (window_videoOut_payload_frame_line_pixel_2_2_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_2_2_15        (window_videoOut_payload_frame_line_pixel_2_2_15[7:0]                    ), //i
    .io_input_payload_frame_line_endOfLine           (window_videoOut_payload_frame_line_endOfLine                            ), //i
    .io_input_payload_frame_endOfFrame               (window_videoOut_payload_frame_endOfFrame                                ), //i
    .io_input_payload_endOfPack                      (window_videoOut_payload_endOfPack                                       ), //i
    .io_outputs_0_valid                              (window_videoOut_fork_io_outputs_0_valid                                 ), //o
    .io_outputs_0_ready                              (unit_0_inputs_ready                                                     ), //i
    .io_outputs_0_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_0_payload_frame_line_endOfLine          ), //o
    .io_outputs_0_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_0_payload_frame_endOfFrame              ), //o
    .io_outputs_0_payload_endOfPack                  (window_videoOut_fork_io_outputs_0_payload_endOfPack                     ), //o
    .io_outputs_1_valid                              (window_videoOut_fork_io_outputs_1_valid                                 ), //o
    .io_outputs_1_ready                              (unit_1_inputs_ready                                                     ), //i
    .io_outputs_1_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_1_payload_frame_line_endOfLine          ), //o
    .io_outputs_1_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_1_payload_frame_endOfFrame              ), //o
    .io_outputs_1_payload_endOfPack                  (window_videoOut_fork_io_outputs_1_payload_endOfPack                     ), //o
    .io_outputs_2_valid                              (window_videoOut_fork_io_outputs_2_valid                                 ), //o
    .io_outputs_2_ready                              (unit_2_inputs_ready                                                     ), //i
    .io_outputs_2_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_2_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_2_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_2_payload_frame_line_endOfLine          ), //o
    .io_outputs_2_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_2_payload_frame_endOfFrame              ), //o
    .io_outputs_2_payload_endOfPack                  (window_videoOut_fork_io_outputs_2_payload_endOfPack                     ), //o
    .io_outputs_3_valid                              (window_videoOut_fork_io_outputs_3_valid                                 ), //o
    .io_outputs_3_ready                              (unit_3_inputs_ready                                                     ), //i
    .io_outputs_3_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_3_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_3_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_3_payload_frame_line_endOfLine          ), //o
    .io_outputs_3_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_3_payload_frame_endOfFrame              ), //o
    .io_outputs_3_payload_endOfPack                  (window_videoOut_fork_io_outputs_3_payload_endOfPack                     ), //o
    .io_outputs_4_valid                              (window_videoOut_fork_io_outputs_4_valid                                 ), //o
    .io_outputs_4_ready                              (unit_4_inputs_ready                                                     ), //i
    .io_outputs_4_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_4_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_4_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_4_payload_frame_line_endOfLine          ), //o
    .io_outputs_4_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_4_payload_frame_endOfFrame              ), //o
    .io_outputs_4_payload_endOfPack                  (window_videoOut_fork_io_outputs_4_payload_endOfPack                     ), //o
    .io_outputs_5_valid                              (window_videoOut_fork_io_outputs_5_valid                                 ), //o
    .io_outputs_5_ready                              (unit_5_inputs_ready                                                     ), //i
    .io_outputs_5_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_5_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_5_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_5_payload_frame_line_endOfLine          ), //o
    .io_outputs_5_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_5_payload_frame_endOfFrame              ), //o
    .io_outputs_5_payload_endOfPack                  (window_videoOut_fork_io_outputs_5_payload_endOfPack                     ), //o
    .io_outputs_6_valid                              (window_videoOut_fork_io_outputs_6_valid                                 ), //o
    .io_outputs_6_ready                              (unit_6_inputs_ready                                                     ), //i
    .io_outputs_6_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_6_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_6_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_6_payload_frame_line_endOfLine          ), //o
    .io_outputs_6_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_6_payload_frame_endOfFrame              ), //o
    .io_outputs_6_payload_endOfPack                  (window_videoOut_fork_io_outputs_6_payload_endOfPack                     ), //o
    .io_outputs_7_valid                              (window_videoOut_fork_io_outputs_7_valid                                 ), //o
    .io_outputs_7_ready                              (unit_7_inputs_ready                                                     ), //i
    .io_outputs_7_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_0[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_1[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_2[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_3[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_4[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_5[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_6[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_7[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_8[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_9[7:0]   ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_10[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_11[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_12[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_13[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_14[7:0]  ), //o
    .io_outputs_7_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_15[7:0]  ), //o
    .io_outputs_7_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_7_payload_frame_line_endOfLine          ), //o
    .io_outputs_7_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_7_payload_frame_endOfFrame              ), //o
    .io_outputs_7_payload_endOfPack                  (window_videoOut_fork_io_outputs_7_payload_endOfPack                     ), //o
    .clk                                             (clk                                                                     ), //i
    .reset                                           (reset                                                                   )  //i
  );
  PecaUnit unit_0 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_0_valid                                 ), //i
    .inputs_ready                              (unit_0_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_0_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_0_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_0_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_0_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_0_pop_valid                                                  ), //i
    .weights_ready                             (unit_0_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_0_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_0_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_0_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_0_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_0_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_0_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_0_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_0_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_0_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_0_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_0_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_0_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_0_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_0_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_0_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_0_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_0_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_0_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_0_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_0_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_0_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_0_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_0_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_0_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_0_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_0_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_0_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_0_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_0_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_0_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_0_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_0_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_0_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_0_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_0_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_0_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_0_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_0_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_0_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_0_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_0_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_0_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_0_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_0_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_0_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_0_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_0_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_0_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_0_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_0_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_0_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_0_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_0_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_0_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_0_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_0_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_0_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_0_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_0_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_0_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_0_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_0_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_0_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_0_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_0_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_0_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_0_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_0_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_0_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_0_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_0_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_0_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_0_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_0_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_0_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_0_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_0_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_0_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_0_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_0_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_0_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_0_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_0_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_0_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_0_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_0_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_0_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_0_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_0_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_0_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_0_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_0_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_0_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_0_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_0_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_0_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_0_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_0_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_0_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_0_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_0_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_0_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_0_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_0_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_0_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_0_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_0_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_0_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_0_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_0_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_0_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_0_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_0_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_0_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_0_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_0_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_0_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_0_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_0_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_0_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_0_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_0_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_0_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_0_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_0_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_0_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_0_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_0_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_0_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_0_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_0_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_0_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_0_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_0_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_0_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_0_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_0_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_0_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_0_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_0_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_0_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_0_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_0_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_0_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_0_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_0_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_0_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_0_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_0_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_0_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_0_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_0_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_0_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_0_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_0_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_0_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_0_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_0_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_0_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_0_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_0_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_0_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_0_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_0_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_0_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_0_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_0_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_0_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_0_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_0_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_0_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_0_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_0_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_0_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_0_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_0_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_0_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_0_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_0_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_0_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_0_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_0_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_0_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_0_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_0_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_0_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_0_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_0_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_0_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_0_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_0_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_0_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_0_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_0_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_0_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_0_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_0_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_0_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_0_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_0_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_0_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_0_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_0_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_0_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_0_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_0_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_0_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_0_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_0_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_0_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_0_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_0_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_0_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_0_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_0_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_0_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_0_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_0_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_0_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_0_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_0_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_0_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_0_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_0_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_0_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_0_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_0_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_0_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_0_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_0_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_0_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_0_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_0_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_0_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_0_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_0_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_0_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_0_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_0_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_0_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_0_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_0_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_0_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_0_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_0_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_0_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_0_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_0_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_0_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_0_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_0_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_0_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_0_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_0_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_0_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_0_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_0_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_0_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_0_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_0_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_0_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_0_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_0_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_0_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_0_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_0_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_0_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_0_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_0_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_0_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_0_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_0_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_0_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_0_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_0_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_0_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_0_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_0_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_0_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_0_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_0_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_0_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_0_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_0_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_0_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_0_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_0_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_0_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_0_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_0_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_0_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_0_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_0_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_0_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_0_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_1 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_1_valid                                 ), //i
    .inputs_ready                              (unit_1_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_1_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_1_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_1_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_1_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_1_pop_valid                                                  ), //i
    .weights_ready                             (unit_1_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_1_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_1_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_1_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_1_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_1_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_1_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_1_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_1_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_1_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_1_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_1_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_1_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_1_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_1_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_1_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_1_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_1_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_1_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_1_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_1_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_1_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_1_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_1_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_1_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_1_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_1_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_1_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_1_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_1_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_1_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_1_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_1_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_1_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_1_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_1_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_1_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_1_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_1_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_1_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_1_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_1_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_1_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_1_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_1_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_1_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_1_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_1_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_1_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_1_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_1_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_1_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_1_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_1_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_1_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_1_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_1_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_1_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_1_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_1_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_1_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_1_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_1_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_1_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_1_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_1_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_1_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_1_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_1_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_1_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_1_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_1_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_1_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_1_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_1_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_1_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_1_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_1_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_1_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_1_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_1_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_1_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_1_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_1_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_1_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_1_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_1_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_1_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_1_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_1_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_1_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_1_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_1_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_1_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_1_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_1_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_1_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_1_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_1_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_1_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_1_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_1_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_1_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_1_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_1_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_1_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_1_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_1_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_1_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_1_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_1_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_1_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_1_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_1_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_1_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_1_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_1_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_1_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_1_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_1_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_1_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_1_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_1_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_1_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_1_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_1_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_1_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_1_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_1_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_1_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_1_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_1_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_1_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_1_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_1_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_1_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_1_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_1_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_1_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_1_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_1_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_1_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_1_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_1_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_1_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_1_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_1_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_1_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_1_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_1_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_1_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_1_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_1_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_1_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_1_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_1_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_1_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_1_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_1_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_1_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_1_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_1_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_1_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_1_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_1_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_1_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_1_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_1_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_1_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_1_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_1_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_1_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_1_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_1_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_1_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_1_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_1_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_1_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_1_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_1_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_1_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_1_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_1_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_1_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_1_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_1_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_1_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_1_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_1_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_1_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_1_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_1_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_1_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_1_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_1_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_1_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_1_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_1_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_1_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_1_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_1_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_1_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_1_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_1_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_1_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_1_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_1_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_1_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_1_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_1_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_1_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_1_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_1_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_1_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_1_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_1_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_1_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_1_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_1_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_1_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_1_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_1_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_1_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_1_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_1_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_1_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_1_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_1_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_1_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_1_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_1_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_1_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_1_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_1_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_1_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_1_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_1_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_1_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_1_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_1_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_1_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_1_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_1_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_1_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_1_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_1_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_1_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_1_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_1_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_1_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_1_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_1_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_1_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_1_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_1_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_1_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_1_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_1_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_1_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_1_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_1_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_1_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_1_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_1_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_1_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_1_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_1_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_1_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_1_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_1_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_1_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_1_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_1_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_1_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_1_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_1_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_1_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_1_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_1_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_1_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_1_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_1_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_1_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_1_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_1_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_1_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_1_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_1_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_1_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_1_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_1_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_1_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_1_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_1_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_1_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_1_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_2 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_2_valid                                 ), //i
    .inputs_ready                              (unit_2_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_2_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_2_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_2_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_2_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_2_pop_valid                                                  ), //i
    .weights_ready                             (unit_2_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_2_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_2_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_2_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_2_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_2_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_2_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_2_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_2_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_2_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_2_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_2_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_2_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_2_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_2_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_2_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_2_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_2_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_2_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_2_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_2_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_2_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_2_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_2_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_2_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_2_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_2_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_2_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_2_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_2_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_2_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_2_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_2_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_2_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_2_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_2_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_2_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_2_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_2_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_2_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_2_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_2_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_2_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_2_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_2_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_2_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_2_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_2_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_2_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_2_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_2_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_2_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_2_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_2_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_2_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_2_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_2_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_2_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_2_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_2_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_2_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_2_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_2_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_2_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_2_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_2_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_2_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_2_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_2_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_2_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_2_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_2_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_2_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_2_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_2_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_2_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_2_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_2_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_2_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_2_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_2_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_2_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_2_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_2_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_2_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_2_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_2_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_2_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_2_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_2_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_2_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_2_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_2_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_2_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_2_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_2_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_2_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_2_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_2_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_2_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_2_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_2_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_2_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_2_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_2_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_2_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_2_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_2_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_2_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_2_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_2_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_2_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_2_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_2_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_2_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_2_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_2_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_2_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_2_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_2_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_2_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_2_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_2_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_2_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_2_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_2_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_2_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_2_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_2_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_2_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_2_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_2_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_2_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_2_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_2_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_2_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_2_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_2_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_2_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_2_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_2_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_2_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_2_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_2_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_2_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_2_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_2_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_2_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_2_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_2_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_2_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_2_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_2_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_2_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_2_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_2_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_2_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_2_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_2_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_2_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_2_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_2_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_2_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_2_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_2_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_2_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_2_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_2_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_2_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_2_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_2_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_2_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_2_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_2_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_2_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_2_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_2_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_2_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_2_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_2_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_2_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_2_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_2_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_2_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_2_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_2_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_2_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_2_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_2_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_2_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_2_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_2_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_2_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_2_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_2_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_2_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_2_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_2_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_2_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_2_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_2_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_2_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_2_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_2_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_2_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_2_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_2_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_2_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_2_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_2_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_2_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_2_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_2_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_2_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_2_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_2_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_2_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_2_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_2_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_2_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_2_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_2_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_2_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_2_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_2_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_2_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_2_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_2_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_2_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_2_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_2_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_2_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_2_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_2_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_2_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_2_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_2_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_2_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_2_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_2_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_2_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_2_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_2_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_2_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_2_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_2_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_2_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_2_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_2_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_2_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_2_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_2_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_2_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_2_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_2_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_2_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_2_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_2_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_2_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_2_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_2_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_2_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_2_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_2_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_2_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_2_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_2_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_2_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_2_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_2_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_2_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_2_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_2_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_2_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_2_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_2_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_2_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_2_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_2_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_2_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_2_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_2_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_2_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_2_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_2_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_2_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_2_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_2_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_2_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_2_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_2_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_2_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_2_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_2_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_2_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_2_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_3 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_3_valid                                 ), //i
    .inputs_ready                              (unit_3_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_3_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_3_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_3_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_3_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_3_pop_valid                                                  ), //i
    .weights_ready                             (unit_3_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_3_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_3_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_3_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_3_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_3_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_3_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_3_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_3_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_3_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_3_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_3_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_3_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_3_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_3_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_3_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_3_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_3_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_3_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_3_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_3_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_3_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_3_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_3_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_3_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_3_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_3_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_3_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_3_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_3_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_3_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_3_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_3_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_3_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_3_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_3_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_3_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_3_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_3_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_3_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_3_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_3_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_3_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_3_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_3_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_3_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_3_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_3_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_3_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_3_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_3_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_3_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_3_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_3_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_3_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_3_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_3_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_3_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_3_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_3_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_3_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_3_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_3_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_3_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_3_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_3_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_3_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_3_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_3_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_3_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_3_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_3_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_3_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_3_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_3_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_3_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_3_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_3_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_3_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_3_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_3_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_3_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_3_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_3_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_3_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_3_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_3_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_3_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_3_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_3_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_3_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_3_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_3_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_3_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_3_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_3_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_3_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_3_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_3_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_3_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_3_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_3_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_3_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_3_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_3_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_3_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_3_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_3_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_3_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_3_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_3_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_3_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_3_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_3_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_3_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_3_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_3_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_3_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_3_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_3_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_3_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_3_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_3_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_3_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_3_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_3_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_3_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_3_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_3_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_3_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_3_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_3_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_3_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_3_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_3_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_3_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_3_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_3_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_3_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_3_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_3_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_3_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_3_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_3_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_3_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_3_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_3_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_3_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_3_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_3_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_3_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_3_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_3_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_3_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_3_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_3_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_3_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_3_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_3_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_3_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_3_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_3_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_3_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_3_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_3_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_3_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_3_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_3_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_3_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_3_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_3_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_3_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_3_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_3_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_3_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_3_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_3_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_3_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_3_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_3_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_3_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_3_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_3_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_3_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_3_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_3_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_3_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_3_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_3_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_3_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_3_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_3_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_3_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_3_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_3_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_3_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_3_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_3_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_3_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_3_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_3_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_3_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_3_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_3_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_3_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_3_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_3_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_3_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_3_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_3_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_3_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_3_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_3_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_3_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_3_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_3_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_3_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_3_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_3_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_3_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_3_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_3_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_3_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_3_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_3_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_3_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_3_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_3_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_3_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_3_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_3_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_3_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_3_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_3_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_3_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_3_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_3_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_3_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_3_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_3_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_3_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_3_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_3_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_3_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_3_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_3_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_3_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_3_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_3_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_3_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_3_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_3_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_3_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_3_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_3_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_3_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_3_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_3_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_3_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_3_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_3_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_3_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_3_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_3_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_3_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_3_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_3_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_3_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_3_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_3_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_3_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_3_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_3_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_3_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_3_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_3_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_3_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_3_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_3_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_3_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_3_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_3_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_3_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_3_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_3_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_3_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_3_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_3_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_3_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_3_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_3_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_3_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_3_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_3_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_3_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_3_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_4 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_4_valid                                 ), //i
    .inputs_ready                              (unit_4_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_4_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_4_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_4_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_4_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_4_pop_valid                                                  ), //i
    .weights_ready                             (unit_4_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_4_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_4_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_4_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_4_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_4_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_4_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_4_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_4_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_4_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_4_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_4_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_4_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_4_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_4_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_4_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_4_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_4_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_4_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_4_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_4_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_4_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_4_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_4_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_4_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_4_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_4_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_4_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_4_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_4_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_4_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_4_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_4_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_4_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_4_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_4_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_4_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_4_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_4_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_4_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_4_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_4_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_4_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_4_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_4_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_4_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_4_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_4_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_4_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_4_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_4_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_4_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_4_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_4_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_4_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_4_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_4_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_4_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_4_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_4_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_4_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_4_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_4_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_4_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_4_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_4_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_4_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_4_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_4_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_4_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_4_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_4_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_4_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_4_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_4_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_4_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_4_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_4_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_4_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_4_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_4_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_4_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_4_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_4_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_4_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_4_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_4_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_4_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_4_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_4_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_4_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_4_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_4_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_4_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_4_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_4_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_4_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_4_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_4_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_4_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_4_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_4_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_4_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_4_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_4_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_4_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_4_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_4_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_4_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_4_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_4_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_4_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_4_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_4_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_4_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_4_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_4_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_4_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_4_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_4_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_4_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_4_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_4_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_4_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_4_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_4_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_4_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_4_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_4_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_4_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_4_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_4_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_4_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_4_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_4_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_4_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_4_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_4_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_4_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_4_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_4_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_4_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_4_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_4_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_4_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_4_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_4_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_4_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_4_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_4_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_4_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_4_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_4_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_4_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_4_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_4_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_4_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_4_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_4_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_4_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_4_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_4_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_4_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_4_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_4_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_4_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_4_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_4_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_4_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_4_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_4_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_4_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_4_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_4_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_4_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_4_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_4_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_4_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_4_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_4_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_4_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_4_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_4_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_4_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_4_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_4_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_4_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_4_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_4_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_4_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_4_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_4_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_4_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_4_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_4_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_4_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_4_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_4_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_4_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_4_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_4_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_4_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_4_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_4_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_4_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_4_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_4_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_4_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_4_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_4_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_4_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_4_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_4_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_4_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_4_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_4_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_4_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_4_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_4_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_4_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_4_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_4_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_4_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_4_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_4_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_4_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_4_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_4_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_4_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_4_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_4_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_4_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_4_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_4_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_4_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_4_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_4_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_4_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_4_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_4_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_4_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_4_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_4_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_4_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_4_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_4_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_4_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_4_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_4_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_4_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_4_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_4_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_4_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_4_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_4_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_4_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_4_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_4_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_4_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_4_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_4_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_4_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_4_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_4_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_4_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_4_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_4_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_4_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_4_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_4_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_4_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_4_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_4_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_4_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_4_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_4_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_4_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_4_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_4_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_4_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_4_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_4_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_4_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_4_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_4_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_4_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_4_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_4_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_4_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_4_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_4_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_4_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_4_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_4_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_4_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_4_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_5 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_5_valid                                 ), //i
    .inputs_ready                              (unit_5_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_5_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_5_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_5_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_5_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_5_pop_valid                                                  ), //i
    .weights_ready                             (unit_5_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_5_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_5_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_5_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_5_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_5_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_5_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_5_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_5_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_5_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_5_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_5_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_5_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_5_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_5_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_5_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_5_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_5_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_5_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_5_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_5_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_5_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_5_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_5_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_5_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_5_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_5_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_5_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_5_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_5_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_5_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_5_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_5_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_5_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_5_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_5_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_5_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_5_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_5_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_5_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_5_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_5_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_5_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_5_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_5_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_5_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_5_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_5_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_5_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_5_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_5_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_5_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_5_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_5_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_5_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_5_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_5_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_5_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_5_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_5_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_5_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_5_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_5_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_5_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_5_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_5_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_5_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_5_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_5_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_5_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_5_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_5_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_5_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_5_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_5_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_5_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_5_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_5_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_5_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_5_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_5_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_5_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_5_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_5_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_5_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_5_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_5_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_5_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_5_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_5_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_5_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_5_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_5_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_5_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_5_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_5_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_5_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_5_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_5_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_5_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_5_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_5_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_5_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_5_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_5_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_5_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_5_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_5_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_5_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_5_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_5_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_5_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_5_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_5_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_5_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_5_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_5_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_5_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_5_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_5_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_5_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_5_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_5_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_5_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_5_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_5_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_5_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_5_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_5_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_5_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_5_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_5_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_5_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_5_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_5_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_5_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_5_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_5_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_5_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_5_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_5_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_5_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_5_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_5_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_5_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_5_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_5_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_5_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_5_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_5_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_5_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_5_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_5_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_5_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_5_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_5_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_5_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_5_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_5_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_5_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_5_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_5_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_5_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_5_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_5_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_5_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_5_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_5_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_5_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_5_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_5_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_5_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_5_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_5_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_5_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_5_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_5_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_5_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_5_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_5_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_5_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_5_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_5_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_5_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_5_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_5_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_5_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_5_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_5_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_5_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_5_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_5_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_5_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_5_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_5_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_5_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_5_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_5_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_5_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_5_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_5_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_5_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_5_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_5_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_5_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_5_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_5_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_5_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_5_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_5_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_5_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_5_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_5_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_5_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_5_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_5_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_5_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_5_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_5_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_5_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_5_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_5_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_5_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_5_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_5_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_5_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_5_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_5_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_5_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_5_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_5_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_5_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_5_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_5_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_5_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_5_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_5_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_5_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_5_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_5_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_5_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_5_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_5_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_5_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_5_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_5_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_5_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_5_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_5_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_5_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_5_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_5_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_5_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_5_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_5_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_5_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_5_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_5_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_5_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_5_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_5_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_5_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_5_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_5_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_5_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_5_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_5_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_5_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_5_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_5_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_5_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_5_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_5_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_5_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_5_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_5_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_5_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_5_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_5_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_5_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_5_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_5_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_5_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_5_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_5_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_5_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_5_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_5_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_5_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_5_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_5_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_5_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_5_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_5_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_5_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_5_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_6 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_6_valid                                 ), //i
    .inputs_ready                              (unit_6_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_6_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_6_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_6_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_6_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_6_pop_valid                                                  ), //i
    .weights_ready                             (unit_6_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_6_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_6_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_6_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_6_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_6_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_6_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_6_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_6_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_6_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_6_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_6_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_6_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_6_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_6_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_6_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_6_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_6_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_6_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_6_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_6_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_6_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_6_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_6_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_6_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_6_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_6_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_6_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_6_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_6_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_6_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_6_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_6_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_6_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_6_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_6_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_6_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_6_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_6_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_6_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_6_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_6_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_6_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_6_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_6_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_6_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_6_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_6_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_6_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_6_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_6_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_6_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_6_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_6_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_6_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_6_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_6_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_6_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_6_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_6_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_6_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_6_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_6_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_6_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_6_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_6_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_6_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_6_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_6_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_6_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_6_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_6_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_6_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_6_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_6_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_6_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_6_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_6_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_6_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_6_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_6_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_6_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_6_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_6_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_6_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_6_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_6_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_6_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_6_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_6_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_6_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_6_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_6_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_6_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_6_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_6_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_6_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_6_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_6_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_6_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_6_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_6_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_6_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_6_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_6_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_6_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_6_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_6_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_6_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_6_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_6_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_6_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_6_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_6_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_6_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_6_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_6_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_6_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_6_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_6_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_6_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_6_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_6_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_6_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_6_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_6_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_6_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_6_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_6_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_6_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_6_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_6_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_6_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_6_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_6_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_6_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_6_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_6_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_6_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_6_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_6_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_6_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_6_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_6_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_6_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_6_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_6_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_6_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_6_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_6_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_6_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_6_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_6_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_6_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_6_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_6_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_6_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_6_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_6_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_6_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_6_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_6_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_6_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_6_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_6_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_6_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_6_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_6_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_6_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_6_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_6_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_6_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_6_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_6_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_6_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_6_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_6_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_6_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_6_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_6_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_6_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_6_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_6_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_6_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_6_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_6_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_6_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_6_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_6_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_6_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_6_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_6_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_6_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_6_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_6_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_6_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_6_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_6_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_6_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_6_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_6_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_6_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_6_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_6_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_6_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_6_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_6_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_6_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_6_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_6_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_6_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_6_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_6_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_6_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_6_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_6_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_6_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_6_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_6_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_6_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_6_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_6_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_6_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_6_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_6_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_6_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_6_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_6_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_6_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_6_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_6_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_6_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_6_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_6_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_6_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_6_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_6_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_6_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_6_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_6_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_6_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_6_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_6_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_6_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_6_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_6_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_6_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_6_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_6_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_6_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_6_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_6_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_6_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_6_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_6_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_6_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_6_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_6_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_6_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_6_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_6_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_6_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_6_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_6_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_6_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_6_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_6_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_6_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_6_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_6_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_6_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_6_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_6_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_6_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_6_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_6_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_6_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_6_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_6_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_6_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_6_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_6_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_6_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_6_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_6_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_6_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_6_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_6_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_6_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_6_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_6_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_6_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_6_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_6_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_6_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_6_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  PecaUnit unit_7 (
    .numberOfInputFrames                       (numberOfInputFrames[7:0]                                                ), //i
    .numberOfOutputFrames                      (numberOfOutputFrames[7:0]                                               ), //i
    .inputs_valid                              (window_videoOut_fork_io_outputs_7_valid                                 ), //i
    .inputs_ready                              (unit_7_inputs_ready                                                     ), //o
    .inputs_payload_frame_line_pixel_0_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_0_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_0_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_0_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_1_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_1_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_1_2_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_0_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_0_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_0_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_1_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_1_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_1_15[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_0     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_0[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_1     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_1[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_2     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_2[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_3     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_3[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_4     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_4[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_5     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_5[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_6     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_6[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_7     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_7[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_8     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_8[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_9     (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_9[7:0]   ), //i
    .inputs_payload_frame_line_pixel_2_2_10    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_10[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_11    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_11[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_12    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_12[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_13    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_13[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_14    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_14[7:0]  ), //i
    .inputs_payload_frame_line_pixel_2_2_15    (window_videoOut_fork_io_outputs_7_payload_frame_line_pixel_2_2_15[7:0]  ), //i
    .inputs_payload_frame_line_endOfLine       (window_videoOut_fork_io_outputs_7_payload_frame_line_endOfLine          ), //i
    .inputs_payload_frame_endOfFrame           (window_videoOut_fork_io_outputs_7_payload_frame_endOfFrame              ), //i
    .inputs_payload_endOfPack                  (window_videoOut_fork_io_outputs_7_payload_endOfPack                     ), //i
    .weights_valid                             (weightFifo_7_pop_valid                                                  ), //i
    .weights_ready                             (unit_7_weights_ready                                                    ), //o
    .weights_payload_0_0_0_0                   (weightFifo_7_pop_payload_0_0_0_0[7:0]                                   ), //i
    .weights_payload_0_0_0_1                   (weightFifo_7_pop_payload_0_0_0_1[7:0]                                   ), //i
    .weights_payload_0_0_0_2                   (weightFifo_7_pop_payload_0_0_0_2[7:0]                                   ), //i
    .weights_payload_0_0_0_3                   (weightFifo_7_pop_payload_0_0_0_3[7:0]                                   ), //i
    .weights_payload_0_0_0_4                   (weightFifo_7_pop_payload_0_0_0_4[7:0]                                   ), //i
    .weights_payload_0_0_0_5                   (weightFifo_7_pop_payload_0_0_0_5[7:0]                                   ), //i
    .weights_payload_0_0_0_6                   (weightFifo_7_pop_payload_0_0_0_6[7:0]                                   ), //i
    .weights_payload_0_0_0_7                   (weightFifo_7_pop_payload_0_0_0_7[7:0]                                   ), //i
    .weights_payload_0_0_0_8                   (weightFifo_7_pop_payload_0_0_0_8[7:0]                                   ), //i
    .weights_payload_0_0_0_9                   (weightFifo_7_pop_payload_0_0_0_9[7:0]                                   ), //i
    .weights_payload_0_0_0_10                  (weightFifo_7_pop_payload_0_0_0_10[7:0]                                  ), //i
    .weights_payload_0_0_0_11                  (weightFifo_7_pop_payload_0_0_0_11[7:0]                                  ), //i
    .weights_payload_0_0_0_12                  (weightFifo_7_pop_payload_0_0_0_12[7:0]                                  ), //i
    .weights_payload_0_0_0_13                  (weightFifo_7_pop_payload_0_0_0_13[7:0]                                  ), //i
    .weights_payload_0_0_0_14                  (weightFifo_7_pop_payload_0_0_0_14[7:0]                                  ), //i
    .weights_payload_0_0_0_15                  (weightFifo_7_pop_payload_0_0_0_15[7:0]                                  ), //i
    .weights_payload_0_0_1_0                   (weightFifo_7_pop_payload_0_0_1_0[7:0]                                   ), //i
    .weights_payload_0_0_1_1                   (weightFifo_7_pop_payload_0_0_1_1[7:0]                                   ), //i
    .weights_payload_0_0_1_2                   (weightFifo_7_pop_payload_0_0_1_2[7:0]                                   ), //i
    .weights_payload_0_0_1_3                   (weightFifo_7_pop_payload_0_0_1_3[7:0]                                   ), //i
    .weights_payload_0_0_1_4                   (weightFifo_7_pop_payload_0_0_1_4[7:0]                                   ), //i
    .weights_payload_0_0_1_5                   (weightFifo_7_pop_payload_0_0_1_5[7:0]                                   ), //i
    .weights_payload_0_0_1_6                   (weightFifo_7_pop_payload_0_0_1_6[7:0]                                   ), //i
    .weights_payload_0_0_1_7                   (weightFifo_7_pop_payload_0_0_1_7[7:0]                                   ), //i
    .weights_payload_0_0_1_8                   (weightFifo_7_pop_payload_0_0_1_8[7:0]                                   ), //i
    .weights_payload_0_0_1_9                   (weightFifo_7_pop_payload_0_0_1_9[7:0]                                   ), //i
    .weights_payload_0_0_1_10                  (weightFifo_7_pop_payload_0_0_1_10[7:0]                                  ), //i
    .weights_payload_0_0_1_11                  (weightFifo_7_pop_payload_0_0_1_11[7:0]                                  ), //i
    .weights_payload_0_0_1_12                  (weightFifo_7_pop_payload_0_0_1_12[7:0]                                  ), //i
    .weights_payload_0_0_1_13                  (weightFifo_7_pop_payload_0_0_1_13[7:0]                                  ), //i
    .weights_payload_0_0_1_14                  (weightFifo_7_pop_payload_0_0_1_14[7:0]                                  ), //i
    .weights_payload_0_0_1_15                  (weightFifo_7_pop_payload_0_0_1_15[7:0]                                  ), //i
    .weights_payload_0_0_2_0                   (weightFifo_7_pop_payload_0_0_2_0[7:0]                                   ), //i
    .weights_payload_0_0_2_1                   (weightFifo_7_pop_payload_0_0_2_1[7:0]                                   ), //i
    .weights_payload_0_0_2_2                   (weightFifo_7_pop_payload_0_0_2_2[7:0]                                   ), //i
    .weights_payload_0_0_2_3                   (weightFifo_7_pop_payload_0_0_2_3[7:0]                                   ), //i
    .weights_payload_0_0_2_4                   (weightFifo_7_pop_payload_0_0_2_4[7:0]                                   ), //i
    .weights_payload_0_0_2_5                   (weightFifo_7_pop_payload_0_0_2_5[7:0]                                   ), //i
    .weights_payload_0_0_2_6                   (weightFifo_7_pop_payload_0_0_2_6[7:0]                                   ), //i
    .weights_payload_0_0_2_7                   (weightFifo_7_pop_payload_0_0_2_7[7:0]                                   ), //i
    .weights_payload_0_0_2_8                   (weightFifo_7_pop_payload_0_0_2_8[7:0]                                   ), //i
    .weights_payload_0_0_2_9                   (weightFifo_7_pop_payload_0_0_2_9[7:0]                                   ), //i
    .weights_payload_0_0_2_10                  (weightFifo_7_pop_payload_0_0_2_10[7:0]                                  ), //i
    .weights_payload_0_0_2_11                  (weightFifo_7_pop_payload_0_0_2_11[7:0]                                  ), //i
    .weights_payload_0_0_2_12                  (weightFifo_7_pop_payload_0_0_2_12[7:0]                                  ), //i
    .weights_payload_0_0_2_13                  (weightFifo_7_pop_payload_0_0_2_13[7:0]                                  ), //i
    .weights_payload_0_0_2_14                  (weightFifo_7_pop_payload_0_0_2_14[7:0]                                  ), //i
    .weights_payload_0_0_2_15                  (weightFifo_7_pop_payload_0_0_2_15[7:0]                                  ), //i
    .weights_payload_0_1_0_0                   (weightFifo_7_pop_payload_0_1_0_0[7:0]                                   ), //i
    .weights_payload_0_1_0_1                   (weightFifo_7_pop_payload_0_1_0_1[7:0]                                   ), //i
    .weights_payload_0_1_0_2                   (weightFifo_7_pop_payload_0_1_0_2[7:0]                                   ), //i
    .weights_payload_0_1_0_3                   (weightFifo_7_pop_payload_0_1_0_3[7:0]                                   ), //i
    .weights_payload_0_1_0_4                   (weightFifo_7_pop_payload_0_1_0_4[7:0]                                   ), //i
    .weights_payload_0_1_0_5                   (weightFifo_7_pop_payload_0_1_0_5[7:0]                                   ), //i
    .weights_payload_0_1_0_6                   (weightFifo_7_pop_payload_0_1_0_6[7:0]                                   ), //i
    .weights_payload_0_1_0_7                   (weightFifo_7_pop_payload_0_1_0_7[7:0]                                   ), //i
    .weights_payload_0_1_0_8                   (weightFifo_7_pop_payload_0_1_0_8[7:0]                                   ), //i
    .weights_payload_0_1_0_9                   (weightFifo_7_pop_payload_0_1_0_9[7:0]                                   ), //i
    .weights_payload_0_1_0_10                  (weightFifo_7_pop_payload_0_1_0_10[7:0]                                  ), //i
    .weights_payload_0_1_0_11                  (weightFifo_7_pop_payload_0_1_0_11[7:0]                                  ), //i
    .weights_payload_0_1_0_12                  (weightFifo_7_pop_payload_0_1_0_12[7:0]                                  ), //i
    .weights_payload_0_1_0_13                  (weightFifo_7_pop_payload_0_1_0_13[7:0]                                  ), //i
    .weights_payload_0_1_0_14                  (weightFifo_7_pop_payload_0_1_0_14[7:0]                                  ), //i
    .weights_payload_0_1_0_15                  (weightFifo_7_pop_payload_0_1_0_15[7:0]                                  ), //i
    .weights_payload_0_1_1_0                   (weightFifo_7_pop_payload_0_1_1_0[7:0]                                   ), //i
    .weights_payload_0_1_1_1                   (weightFifo_7_pop_payload_0_1_1_1[7:0]                                   ), //i
    .weights_payload_0_1_1_2                   (weightFifo_7_pop_payload_0_1_1_2[7:0]                                   ), //i
    .weights_payload_0_1_1_3                   (weightFifo_7_pop_payload_0_1_1_3[7:0]                                   ), //i
    .weights_payload_0_1_1_4                   (weightFifo_7_pop_payload_0_1_1_4[7:0]                                   ), //i
    .weights_payload_0_1_1_5                   (weightFifo_7_pop_payload_0_1_1_5[7:0]                                   ), //i
    .weights_payload_0_1_1_6                   (weightFifo_7_pop_payload_0_1_1_6[7:0]                                   ), //i
    .weights_payload_0_1_1_7                   (weightFifo_7_pop_payload_0_1_1_7[7:0]                                   ), //i
    .weights_payload_0_1_1_8                   (weightFifo_7_pop_payload_0_1_1_8[7:0]                                   ), //i
    .weights_payload_0_1_1_9                   (weightFifo_7_pop_payload_0_1_1_9[7:0]                                   ), //i
    .weights_payload_0_1_1_10                  (weightFifo_7_pop_payload_0_1_1_10[7:0]                                  ), //i
    .weights_payload_0_1_1_11                  (weightFifo_7_pop_payload_0_1_1_11[7:0]                                  ), //i
    .weights_payload_0_1_1_12                  (weightFifo_7_pop_payload_0_1_1_12[7:0]                                  ), //i
    .weights_payload_0_1_1_13                  (weightFifo_7_pop_payload_0_1_1_13[7:0]                                  ), //i
    .weights_payload_0_1_1_14                  (weightFifo_7_pop_payload_0_1_1_14[7:0]                                  ), //i
    .weights_payload_0_1_1_15                  (weightFifo_7_pop_payload_0_1_1_15[7:0]                                  ), //i
    .weights_payload_0_1_2_0                   (weightFifo_7_pop_payload_0_1_2_0[7:0]                                   ), //i
    .weights_payload_0_1_2_1                   (weightFifo_7_pop_payload_0_1_2_1[7:0]                                   ), //i
    .weights_payload_0_1_2_2                   (weightFifo_7_pop_payload_0_1_2_2[7:0]                                   ), //i
    .weights_payload_0_1_2_3                   (weightFifo_7_pop_payload_0_1_2_3[7:0]                                   ), //i
    .weights_payload_0_1_2_4                   (weightFifo_7_pop_payload_0_1_2_4[7:0]                                   ), //i
    .weights_payload_0_1_2_5                   (weightFifo_7_pop_payload_0_1_2_5[7:0]                                   ), //i
    .weights_payload_0_1_2_6                   (weightFifo_7_pop_payload_0_1_2_6[7:0]                                   ), //i
    .weights_payload_0_1_2_7                   (weightFifo_7_pop_payload_0_1_2_7[7:0]                                   ), //i
    .weights_payload_0_1_2_8                   (weightFifo_7_pop_payload_0_1_2_8[7:0]                                   ), //i
    .weights_payload_0_1_2_9                   (weightFifo_7_pop_payload_0_1_2_9[7:0]                                   ), //i
    .weights_payload_0_1_2_10                  (weightFifo_7_pop_payload_0_1_2_10[7:0]                                  ), //i
    .weights_payload_0_1_2_11                  (weightFifo_7_pop_payload_0_1_2_11[7:0]                                  ), //i
    .weights_payload_0_1_2_12                  (weightFifo_7_pop_payload_0_1_2_12[7:0]                                  ), //i
    .weights_payload_0_1_2_13                  (weightFifo_7_pop_payload_0_1_2_13[7:0]                                  ), //i
    .weights_payload_0_1_2_14                  (weightFifo_7_pop_payload_0_1_2_14[7:0]                                  ), //i
    .weights_payload_0_1_2_15                  (weightFifo_7_pop_payload_0_1_2_15[7:0]                                  ), //i
    .weights_payload_0_2_0_0                   (weightFifo_7_pop_payload_0_2_0_0[7:0]                                   ), //i
    .weights_payload_0_2_0_1                   (weightFifo_7_pop_payload_0_2_0_1[7:0]                                   ), //i
    .weights_payload_0_2_0_2                   (weightFifo_7_pop_payload_0_2_0_2[7:0]                                   ), //i
    .weights_payload_0_2_0_3                   (weightFifo_7_pop_payload_0_2_0_3[7:0]                                   ), //i
    .weights_payload_0_2_0_4                   (weightFifo_7_pop_payload_0_2_0_4[7:0]                                   ), //i
    .weights_payload_0_2_0_5                   (weightFifo_7_pop_payload_0_2_0_5[7:0]                                   ), //i
    .weights_payload_0_2_0_6                   (weightFifo_7_pop_payload_0_2_0_6[7:0]                                   ), //i
    .weights_payload_0_2_0_7                   (weightFifo_7_pop_payload_0_2_0_7[7:0]                                   ), //i
    .weights_payload_0_2_0_8                   (weightFifo_7_pop_payload_0_2_0_8[7:0]                                   ), //i
    .weights_payload_0_2_0_9                   (weightFifo_7_pop_payload_0_2_0_9[7:0]                                   ), //i
    .weights_payload_0_2_0_10                  (weightFifo_7_pop_payload_0_2_0_10[7:0]                                  ), //i
    .weights_payload_0_2_0_11                  (weightFifo_7_pop_payload_0_2_0_11[7:0]                                  ), //i
    .weights_payload_0_2_0_12                  (weightFifo_7_pop_payload_0_2_0_12[7:0]                                  ), //i
    .weights_payload_0_2_0_13                  (weightFifo_7_pop_payload_0_2_0_13[7:0]                                  ), //i
    .weights_payload_0_2_0_14                  (weightFifo_7_pop_payload_0_2_0_14[7:0]                                  ), //i
    .weights_payload_0_2_0_15                  (weightFifo_7_pop_payload_0_2_0_15[7:0]                                  ), //i
    .weights_payload_0_2_1_0                   (weightFifo_7_pop_payload_0_2_1_0[7:0]                                   ), //i
    .weights_payload_0_2_1_1                   (weightFifo_7_pop_payload_0_2_1_1[7:0]                                   ), //i
    .weights_payload_0_2_1_2                   (weightFifo_7_pop_payload_0_2_1_2[7:0]                                   ), //i
    .weights_payload_0_2_1_3                   (weightFifo_7_pop_payload_0_2_1_3[7:0]                                   ), //i
    .weights_payload_0_2_1_4                   (weightFifo_7_pop_payload_0_2_1_4[7:0]                                   ), //i
    .weights_payload_0_2_1_5                   (weightFifo_7_pop_payload_0_2_1_5[7:0]                                   ), //i
    .weights_payload_0_2_1_6                   (weightFifo_7_pop_payload_0_2_1_6[7:0]                                   ), //i
    .weights_payload_0_2_1_7                   (weightFifo_7_pop_payload_0_2_1_7[7:0]                                   ), //i
    .weights_payload_0_2_1_8                   (weightFifo_7_pop_payload_0_2_1_8[7:0]                                   ), //i
    .weights_payload_0_2_1_9                   (weightFifo_7_pop_payload_0_2_1_9[7:0]                                   ), //i
    .weights_payload_0_2_1_10                  (weightFifo_7_pop_payload_0_2_1_10[7:0]                                  ), //i
    .weights_payload_0_2_1_11                  (weightFifo_7_pop_payload_0_2_1_11[7:0]                                  ), //i
    .weights_payload_0_2_1_12                  (weightFifo_7_pop_payload_0_2_1_12[7:0]                                  ), //i
    .weights_payload_0_2_1_13                  (weightFifo_7_pop_payload_0_2_1_13[7:0]                                  ), //i
    .weights_payload_0_2_1_14                  (weightFifo_7_pop_payload_0_2_1_14[7:0]                                  ), //i
    .weights_payload_0_2_1_15                  (weightFifo_7_pop_payload_0_2_1_15[7:0]                                  ), //i
    .weights_payload_0_2_2_0                   (weightFifo_7_pop_payload_0_2_2_0[7:0]                                   ), //i
    .weights_payload_0_2_2_1                   (weightFifo_7_pop_payload_0_2_2_1[7:0]                                   ), //i
    .weights_payload_0_2_2_2                   (weightFifo_7_pop_payload_0_2_2_2[7:0]                                   ), //i
    .weights_payload_0_2_2_3                   (weightFifo_7_pop_payload_0_2_2_3[7:0]                                   ), //i
    .weights_payload_0_2_2_4                   (weightFifo_7_pop_payload_0_2_2_4[7:0]                                   ), //i
    .weights_payload_0_2_2_5                   (weightFifo_7_pop_payload_0_2_2_5[7:0]                                   ), //i
    .weights_payload_0_2_2_6                   (weightFifo_7_pop_payload_0_2_2_6[7:0]                                   ), //i
    .weights_payload_0_2_2_7                   (weightFifo_7_pop_payload_0_2_2_7[7:0]                                   ), //i
    .weights_payload_0_2_2_8                   (weightFifo_7_pop_payload_0_2_2_8[7:0]                                   ), //i
    .weights_payload_0_2_2_9                   (weightFifo_7_pop_payload_0_2_2_9[7:0]                                   ), //i
    .weights_payload_0_2_2_10                  (weightFifo_7_pop_payload_0_2_2_10[7:0]                                  ), //i
    .weights_payload_0_2_2_11                  (weightFifo_7_pop_payload_0_2_2_11[7:0]                                  ), //i
    .weights_payload_0_2_2_12                  (weightFifo_7_pop_payload_0_2_2_12[7:0]                                  ), //i
    .weights_payload_0_2_2_13                  (weightFifo_7_pop_payload_0_2_2_13[7:0]                                  ), //i
    .weights_payload_0_2_2_14                  (weightFifo_7_pop_payload_0_2_2_14[7:0]                                  ), //i
    .weights_payload_0_2_2_15                  (weightFifo_7_pop_payload_0_2_2_15[7:0]                                  ), //i
    .weights_payload_1_0_0_0                   (weightFifo_7_pop_payload_1_0_0_0[7:0]                                   ), //i
    .weights_payload_1_0_0_1                   (weightFifo_7_pop_payload_1_0_0_1[7:0]                                   ), //i
    .weights_payload_1_0_0_2                   (weightFifo_7_pop_payload_1_0_0_2[7:0]                                   ), //i
    .weights_payload_1_0_0_3                   (weightFifo_7_pop_payload_1_0_0_3[7:0]                                   ), //i
    .weights_payload_1_0_0_4                   (weightFifo_7_pop_payload_1_0_0_4[7:0]                                   ), //i
    .weights_payload_1_0_0_5                   (weightFifo_7_pop_payload_1_0_0_5[7:0]                                   ), //i
    .weights_payload_1_0_0_6                   (weightFifo_7_pop_payload_1_0_0_6[7:0]                                   ), //i
    .weights_payload_1_0_0_7                   (weightFifo_7_pop_payload_1_0_0_7[7:0]                                   ), //i
    .weights_payload_1_0_0_8                   (weightFifo_7_pop_payload_1_0_0_8[7:0]                                   ), //i
    .weights_payload_1_0_0_9                   (weightFifo_7_pop_payload_1_0_0_9[7:0]                                   ), //i
    .weights_payload_1_0_0_10                  (weightFifo_7_pop_payload_1_0_0_10[7:0]                                  ), //i
    .weights_payload_1_0_0_11                  (weightFifo_7_pop_payload_1_0_0_11[7:0]                                  ), //i
    .weights_payload_1_0_0_12                  (weightFifo_7_pop_payload_1_0_0_12[7:0]                                  ), //i
    .weights_payload_1_0_0_13                  (weightFifo_7_pop_payload_1_0_0_13[7:0]                                  ), //i
    .weights_payload_1_0_0_14                  (weightFifo_7_pop_payload_1_0_0_14[7:0]                                  ), //i
    .weights_payload_1_0_0_15                  (weightFifo_7_pop_payload_1_0_0_15[7:0]                                  ), //i
    .weights_payload_1_0_1_0                   (weightFifo_7_pop_payload_1_0_1_0[7:0]                                   ), //i
    .weights_payload_1_0_1_1                   (weightFifo_7_pop_payload_1_0_1_1[7:0]                                   ), //i
    .weights_payload_1_0_1_2                   (weightFifo_7_pop_payload_1_0_1_2[7:0]                                   ), //i
    .weights_payload_1_0_1_3                   (weightFifo_7_pop_payload_1_0_1_3[7:0]                                   ), //i
    .weights_payload_1_0_1_4                   (weightFifo_7_pop_payload_1_0_1_4[7:0]                                   ), //i
    .weights_payload_1_0_1_5                   (weightFifo_7_pop_payload_1_0_1_5[7:0]                                   ), //i
    .weights_payload_1_0_1_6                   (weightFifo_7_pop_payload_1_0_1_6[7:0]                                   ), //i
    .weights_payload_1_0_1_7                   (weightFifo_7_pop_payload_1_0_1_7[7:0]                                   ), //i
    .weights_payload_1_0_1_8                   (weightFifo_7_pop_payload_1_0_1_8[7:0]                                   ), //i
    .weights_payload_1_0_1_9                   (weightFifo_7_pop_payload_1_0_1_9[7:0]                                   ), //i
    .weights_payload_1_0_1_10                  (weightFifo_7_pop_payload_1_0_1_10[7:0]                                  ), //i
    .weights_payload_1_0_1_11                  (weightFifo_7_pop_payload_1_0_1_11[7:0]                                  ), //i
    .weights_payload_1_0_1_12                  (weightFifo_7_pop_payload_1_0_1_12[7:0]                                  ), //i
    .weights_payload_1_0_1_13                  (weightFifo_7_pop_payload_1_0_1_13[7:0]                                  ), //i
    .weights_payload_1_0_1_14                  (weightFifo_7_pop_payload_1_0_1_14[7:0]                                  ), //i
    .weights_payload_1_0_1_15                  (weightFifo_7_pop_payload_1_0_1_15[7:0]                                  ), //i
    .weights_payload_1_0_2_0                   (weightFifo_7_pop_payload_1_0_2_0[7:0]                                   ), //i
    .weights_payload_1_0_2_1                   (weightFifo_7_pop_payload_1_0_2_1[7:0]                                   ), //i
    .weights_payload_1_0_2_2                   (weightFifo_7_pop_payload_1_0_2_2[7:0]                                   ), //i
    .weights_payload_1_0_2_3                   (weightFifo_7_pop_payload_1_0_2_3[7:0]                                   ), //i
    .weights_payload_1_0_2_4                   (weightFifo_7_pop_payload_1_0_2_4[7:0]                                   ), //i
    .weights_payload_1_0_2_5                   (weightFifo_7_pop_payload_1_0_2_5[7:0]                                   ), //i
    .weights_payload_1_0_2_6                   (weightFifo_7_pop_payload_1_0_2_6[7:0]                                   ), //i
    .weights_payload_1_0_2_7                   (weightFifo_7_pop_payload_1_0_2_7[7:0]                                   ), //i
    .weights_payload_1_0_2_8                   (weightFifo_7_pop_payload_1_0_2_8[7:0]                                   ), //i
    .weights_payload_1_0_2_9                   (weightFifo_7_pop_payload_1_0_2_9[7:0]                                   ), //i
    .weights_payload_1_0_2_10                  (weightFifo_7_pop_payload_1_0_2_10[7:0]                                  ), //i
    .weights_payload_1_0_2_11                  (weightFifo_7_pop_payload_1_0_2_11[7:0]                                  ), //i
    .weights_payload_1_0_2_12                  (weightFifo_7_pop_payload_1_0_2_12[7:0]                                  ), //i
    .weights_payload_1_0_2_13                  (weightFifo_7_pop_payload_1_0_2_13[7:0]                                  ), //i
    .weights_payload_1_0_2_14                  (weightFifo_7_pop_payload_1_0_2_14[7:0]                                  ), //i
    .weights_payload_1_0_2_15                  (weightFifo_7_pop_payload_1_0_2_15[7:0]                                  ), //i
    .weights_payload_1_1_0_0                   (weightFifo_7_pop_payload_1_1_0_0[7:0]                                   ), //i
    .weights_payload_1_1_0_1                   (weightFifo_7_pop_payload_1_1_0_1[7:0]                                   ), //i
    .weights_payload_1_1_0_2                   (weightFifo_7_pop_payload_1_1_0_2[7:0]                                   ), //i
    .weights_payload_1_1_0_3                   (weightFifo_7_pop_payload_1_1_0_3[7:0]                                   ), //i
    .weights_payload_1_1_0_4                   (weightFifo_7_pop_payload_1_1_0_4[7:0]                                   ), //i
    .weights_payload_1_1_0_5                   (weightFifo_7_pop_payload_1_1_0_5[7:0]                                   ), //i
    .weights_payload_1_1_0_6                   (weightFifo_7_pop_payload_1_1_0_6[7:0]                                   ), //i
    .weights_payload_1_1_0_7                   (weightFifo_7_pop_payload_1_1_0_7[7:0]                                   ), //i
    .weights_payload_1_1_0_8                   (weightFifo_7_pop_payload_1_1_0_8[7:0]                                   ), //i
    .weights_payload_1_1_0_9                   (weightFifo_7_pop_payload_1_1_0_9[7:0]                                   ), //i
    .weights_payload_1_1_0_10                  (weightFifo_7_pop_payload_1_1_0_10[7:0]                                  ), //i
    .weights_payload_1_1_0_11                  (weightFifo_7_pop_payload_1_1_0_11[7:0]                                  ), //i
    .weights_payload_1_1_0_12                  (weightFifo_7_pop_payload_1_1_0_12[7:0]                                  ), //i
    .weights_payload_1_1_0_13                  (weightFifo_7_pop_payload_1_1_0_13[7:0]                                  ), //i
    .weights_payload_1_1_0_14                  (weightFifo_7_pop_payload_1_1_0_14[7:0]                                  ), //i
    .weights_payload_1_1_0_15                  (weightFifo_7_pop_payload_1_1_0_15[7:0]                                  ), //i
    .weights_payload_1_1_1_0                   (weightFifo_7_pop_payload_1_1_1_0[7:0]                                   ), //i
    .weights_payload_1_1_1_1                   (weightFifo_7_pop_payload_1_1_1_1[7:0]                                   ), //i
    .weights_payload_1_1_1_2                   (weightFifo_7_pop_payload_1_1_1_2[7:0]                                   ), //i
    .weights_payload_1_1_1_3                   (weightFifo_7_pop_payload_1_1_1_3[7:0]                                   ), //i
    .weights_payload_1_1_1_4                   (weightFifo_7_pop_payload_1_1_1_4[7:0]                                   ), //i
    .weights_payload_1_1_1_5                   (weightFifo_7_pop_payload_1_1_1_5[7:0]                                   ), //i
    .weights_payload_1_1_1_6                   (weightFifo_7_pop_payload_1_1_1_6[7:0]                                   ), //i
    .weights_payload_1_1_1_7                   (weightFifo_7_pop_payload_1_1_1_7[7:0]                                   ), //i
    .weights_payload_1_1_1_8                   (weightFifo_7_pop_payload_1_1_1_8[7:0]                                   ), //i
    .weights_payload_1_1_1_9                   (weightFifo_7_pop_payload_1_1_1_9[7:0]                                   ), //i
    .weights_payload_1_1_1_10                  (weightFifo_7_pop_payload_1_1_1_10[7:0]                                  ), //i
    .weights_payload_1_1_1_11                  (weightFifo_7_pop_payload_1_1_1_11[7:0]                                  ), //i
    .weights_payload_1_1_1_12                  (weightFifo_7_pop_payload_1_1_1_12[7:0]                                  ), //i
    .weights_payload_1_1_1_13                  (weightFifo_7_pop_payload_1_1_1_13[7:0]                                  ), //i
    .weights_payload_1_1_1_14                  (weightFifo_7_pop_payload_1_1_1_14[7:0]                                  ), //i
    .weights_payload_1_1_1_15                  (weightFifo_7_pop_payload_1_1_1_15[7:0]                                  ), //i
    .weights_payload_1_1_2_0                   (weightFifo_7_pop_payload_1_1_2_0[7:0]                                   ), //i
    .weights_payload_1_1_2_1                   (weightFifo_7_pop_payload_1_1_2_1[7:0]                                   ), //i
    .weights_payload_1_1_2_2                   (weightFifo_7_pop_payload_1_1_2_2[7:0]                                   ), //i
    .weights_payload_1_1_2_3                   (weightFifo_7_pop_payload_1_1_2_3[7:0]                                   ), //i
    .weights_payload_1_1_2_4                   (weightFifo_7_pop_payload_1_1_2_4[7:0]                                   ), //i
    .weights_payload_1_1_2_5                   (weightFifo_7_pop_payload_1_1_2_5[7:0]                                   ), //i
    .weights_payload_1_1_2_6                   (weightFifo_7_pop_payload_1_1_2_6[7:0]                                   ), //i
    .weights_payload_1_1_2_7                   (weightFifo_7_pop_payload_1_1_2_7[7:0]                                   ), //i
    .weights_payload_1_1_2_8                   (weightFifo_7_pop_payload_1_1_2_8[7:0]                                   ), //i
    .weights_payload_1_1_2_9                   (weightFifo_7_pop_payload_1_1_2_9[7:0]                                   ), //i
    .weights_payload_1_1_2_10                  (weightFifo_7_pop_payload_1_1_2_10[7:0]                                  ), //i
    .weights_payload_1_1_2_11                  (weightFifo_7_pop_payload_1_1_2_11[7:0]                                  ), //i
    .weights_payload_1_1_2_12                  (weightFifo_7_pop_payload_1_1_2_12[7:0]                                  ), //i
    .weights_payload_1_1_2_13                  (weightFifo_7_pop_payload_1_1_2_13[7:0]                                  ), //i
    .weights_payload_1_1_2_14                  (weightFifo_7_pop_payload_1_1_2_14[7:0]                                  ), //i
    .weights_payload_1_1_2_15                  (weightFifo_7_pop_payload_1_1_2_15[7:0]                                  ), //i
    .weights_payload_1_2_0_0                   (weightFifo_7_pop_payload_1_2_0_0[7:0]                                   ), //i
    .weights_payload_1_2_0_1                   (weightFifo_7_pop_payload_1_2_0_1[7:0]                                   ), //i
    .weights_payload_1_2_0_2                   (weightFifo_7_pop_payload_1_2_0_2[7:0]                                   ), //i
    .weights_payload_1_2_0_3                   (weightFifo_7_pop_payload_1_2_0_3[7:0]                                   ), //i
    .weights_payload_1_2_0_4                   (weightFifo_7_pop_payload_1_2_0_4[7:0]                                   ), //i
    .weights_payload_1_2_0_5                   (weightFifo_7_pop_payload_1_2_0_5[7:0]                                   ), //i
    .weights_payload_1_2_0_6                   (weightFifo_7_pop_payload_1_2_0_6[7:0]                                   ), //i
    .weights_payload_1_2_0_7                   (weightFifo_7_pop_payload_1_2_0_7[7:0]                                   ), //i
    .weights_payload_1_2_0_8                   (weightFifo_7_pop_payload_1_2_0_8[7:0]                                   ), //i
    .weights_payload_1_2_0_9                   (weightFifo_7_pop_payload_1_2_0_9[7:0]                                   ), //i
    .weights_payload_1_2_0_10                  (weightFifo_7_pop_payload_1_2_0_10[7:0]                                  ), //i
    .weights_payload_1_2_0_11                  (weightFifo_7_pop_payload_1_2_0_11[7:0]                                  ), //i
    .weights_payload_1_2_0_12                  (weightFifo_7_pop_payload_1_2_0_12[7:0]                                  ), //i
    .weights_payload_1_2_0_13                  (weightFifo_7_pop_payload_1_2_0_13[7:0]                                  ), //i
    .weights_payload_1_2_0_14                  (weightFifo_7_pop_payload_1_2_0_14[7:0]                                  ), //i
    .weights_payload_1_2_0_15                  (weightFifo_7_pop_payload_1_2_0_15[7:0]                                  ), //i
    .weights_payload_1_2_1_0                   (weightFifo_7_pop_payload_1_2_1_0[7:0]                                   ), //i
    .weights_payload_1_2_1_1                   (weightFifo_7_pop_payload_1_2_1_1[7:0]                                   ), //i
    .weights_payload_1_2_1_2                   (weightFifo_7_pop_payload_1_2_1_2[7:0]                                   ), //i
    .weights_payload_1_2_1_3                   (weightFifo_7_pop_payload_1_2_1_3[7:0]                                   ), //i
    .weights_payload_1_2_1_4                   (weightFifo_7_pop_payload_1_2_1_4[7:0]                                   ), //i
    .weights_payload_1_2_1_5                   (weightFifo_7_pop_payload_1_2_1_5[7:0]                                   ), //i
    .weights_payload_1_2_1_6                   (weightFifo_7_pop_payload_1_2_1_6[7:0]                                   ), //i
    .weights_payload_1_2_1_7                   (weightFifo_7_pop_payload_1_2_1_7[7:0]                                   ), //i
    .weights_payload_1_2_1_8                   (weightFifo_7_pop_payload_1_2_1_8[7:0]                                   ), //i
    .weights_payload_1_2_1_9                   (weightFifo_7_pop_payload_1_2_1_9[7:0]                                   ), //i
    .weights_payload_1_2_1_10                  (weightFifo_7_pop_payload_1_2_1_10[7:0]                                  ), //i
    .weights_payload_1_2_1_11                  (weightFifo_7_pop_payload_1_2_1_11[7:0]                                  ), //i
    .weights_payload_1_2_1_12                  (weightFifo_7_pop_payload_1_2_1_12[7:0]                                  ), //i
    .weights_payload_1_2_1_13                  (weightFifo_7_pop_payload_1_2_1_13[7:0]                                  ), //i
    .weights_payload_1_2_1_14                  (weightFifo_7_pop_payload_1_2_1_14[7:0]                                  ), //i
    .weights_payload_1_2_1_15                  (weightFifo_7_pop_payload_1_2_1_15[7:0]                                  ), //i
    .weights_payload_1_2_2_0                   (weightFifo_7_pop_payload_1_2_2_0[7:0]                                   ), //i
    .weights_payload_1_2_2_1                   (weightFifo_7_pop_payload_1_2_2_1[7:0]                                   ), //i
    .weights_payload_1_2_2_2                   (weightFifo_7_pop_payload_1_2_2_2[7:0]                                   ), //i
    .weights_payload_1_2_2_3                   (weightFifo_7_pop_payload_1_2_2_3[7:0]                                   ), //i
    .weights_payload_1_2_2_4                   (weightFifo_7_pop_payload_1_2_2_4[7:0]                                   ), //i
    .weights_payload_1_2_2_5                   (weightFifo_7_pop_payload_1_2_2_5[7:0]                                   ), //i
    .weights_payload_1_2_2_6                   (weightFifo_7_pop_payload_1_2_2_6[7:0]                                   ), //i
    .weights_payload_1_2_2_7                   (weightFifo_7_pop_payload_1_2_2_7[7:0]                                   ), //i
    .weights_payload_1_2_2_8                   (weightFifo_7_pop_payload_1_2_2_8[7:0]                                   ), //i
    .weights_payload_1_2_2_9                   (weightFifo_7_pop_payload_1_2_2_9[7:0]                                   ), //i
    .weights_payload_1_2_2_10                  (weightFifo_7_pop_payload_1_2_2_10[7:0]                                  ), //i
    .weights_payload_1_2_2_11                  (weightFifo_7_pop_payload_1_2_2_11[7:0]                                  ), //i
    .weights_payload_1_2_2_12                  (weightFifo_7_pop_payload_1_2_2_12[7:0]                                  ), //i
    .weights_payload_1_2_2_13                  (weightFifo_7_pop_payload_1_2_2_13[7:0]                                  ), //i
    .weights_payload_1_2_2_14                  (weightFifo_7_pop_payload_1_2_2_14[7:0]                                  ), //i
    .weights_payload_1_2_2_15                  (weightFifo_7_pop_payload_1_2_2_15[7:0]                                  ), //i
    .outputs_valid                             (unit_7_outputs_valid                                                    ), //o
    .outputs_ready                             (accOutputs_7_ready                                                      ), //i
    .outputs_payload_frame_line_pixel_0        (unit_7_outputs_payload_frame_line_pixel_0[23:0]                         ), //o
    .outputs_payload_frame_line_pixel_1        (unit_7_outputs_payload_frame_line_pixel_1[23:0]                         ), //o
    .outputs_payload_frame_line_endOfLine      (unit_7_outputs_payload_frame_line_endOfLine                             ), //o
    .outputs_payload_frame_endOfFrame          (unit_7_outputs_payload_frame_endOfFrame                                 ), //o
    .outputs_payload_endOfPack                 (unit_7_outputs_payload_endOfPack                                        ), //o
    .clk                                       (clk                                                                     ), //i
    .reset                                     (reset                                                                   )  //i
  );
  VideoPooling pool (
    .videoIn_valid                            (streamDemux_3_io_outputs_1_valid                             ), //i
    .videoIn_ready                            (pool_videoIn_ready                                           ), //o
    .videoIn_payload_frame_line_pixel_0       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_3       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_4       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_5       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_6       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_7       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_8       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_9       (streamDemux_3_io_outputs_1_payload_frame_line_pixel_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_10      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_11      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_12      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_13      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_14      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_15      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_15[7:0]  ), //i
    .videoIn_payload_frame_line_endOfLine     (streamDemux_3_io_outputs_1_payload_frame_line_endOfLine      ), //i
    .videoIn_payload_frame_endOfFrame         (streamDemux_3_io_outputs_1_payload_frame_endOfFrame          ), //i
    .videoIn_payload_endOfPack                (streamDemux_3_io_outputs_1_payload_endOfPack                 ), //i
    .videoOut_valid                           (pool_videoOut_valid                                          ), //o
    .videoOut_ready                           (streamMux_1_io_inputs_1_ready                                ), //i
    .videoOut_payload_frame_line_pixel_0      (pool_videoOut_payload_frame_line_pixel_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1      (pool_videoOut_payload_frame_line_pixel_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2      (pool_videoOut_payload_frame_line_pixel_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_3      (pool_videoOut_payload_frame_line_pixel_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_4      (pool_videoOut_payload_frame_line_pixel_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_5      (pool_videoOut_payload_frame_line_pixel_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_6      (pool_videoOut_payload_frame_line_pixel_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_7      (pool_videoOut_payload_frame_line_pixel_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_8      (pool_videoOut_payload_frame_line_pixel_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_9      (pool_videoOut_payload_frame_line_pixel_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_10     (pool_videoOut_payload_frame_line_pixel_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_11     (pool_videoOut_payload_frame_line_pixel_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_12     (pool_videoOut_payload_frame_line_pixel_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_13     (pool_videoOut_payload_frame_line_pixel_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_14     (pool_videoOut_payload_frame_line_pixel_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_15     (pool_videoOut_payload_frame_line_pixel_15[7:0]               ), //o
    .videoOut_payload_frame_line_endOfLine    (pool_videoOut_payload_frame_line_endOfLine                   ), //o
    .videoOut_payload_frame_endOfFrame        (pool_videoOut_payload_frame_endOfFrame                       ), //o
    .videoOut_payload_endOfPack               (pool_videoOut_payload_endOfPack                              ), //o
    .clk                                      (clk                                                          ), //i
    .reset                                    (reset                                                        )  //i
  );
  LookUpTable table_1 (
    .newTable_valid      (tableAdapted_valid              ), //i
    .newTable_ready      (table_1_newTable_ready          ), //o
    .newTable_payload    (tableAdapted_payload[7:0]       ), //i
    .index_valid         (signalTrim_valid                ), //i
    .index_ready         (table_1_index_ready             ), //o
    .index_payload_0     (signalTrim_payload_0[7:0]       ), //i
    .index_payload_1     (signalTrim_payload_1[7:0]       ), //i
    .index_payload_2     (signalTrim_payload_2[7:0]       ), //i
    .index_payload_3     (signalTrim_payload_3[7:0]       ), //i
    .index_payload_4     (signalTrim_payload_4[7:0]       ), //i
    .index_payload_5     (signalTrim_payload_5[7:0]       ), //i
    .index_payload_6     (signalTrim_payload_6[7:0]       ), //i
    .index_payload_7     (signalTrim_payload_7[7:0]       ), //i
    .index_payload_8     (signalTrim_payload_8[7:0]       ), //i
    .index_payload_9     (signalTrim_payload_9[7:0]       ), //i
    .index_payload_10    (signalTrim_payload_10[7:0]      ), //i
    .index_payload_11    (signalTrim_payload_11[7:0]      ), //i
    .index_payload_12    (signalTrim_payload_12[7:0]      ), //i
    .index_payload_13    (signalTrim_payload_13[7:0]      ), //i
    .index_payload_14    (signalTrim_payload_14[7:0]      ), //i
    .index_payload_15    (signalTrim_payload_15[7:0]      ), //i
    .value_valid         (table_1_value_valid             ), //o
    .value_ready         (table_1_value_transmuted_ready  ), //i
    .value_payload_0     (table_1_value_payload_0[7:0]    ), //o
    .value_payload_1     (table_1_value_payload_1[7:0]    ), //o
    .value_payload_2     (table_1_value_payload_2[7:0]    ), //o
    .value_payload_3     (table_1_value_payload_3[7:0]    ), //o
    .value_payload_4     (table_1_value_payload_4[7:0]    ), //o
    .value_payload_5     (table_1_value_payload_5[7:0]    ), //o
    .value_payload_6     (table_1_value_payload_6[7:0]    ), //o
    .value_payload_7     (table_1_value_payload_7[7:0]    ), //o
    .value_payload_8     (table_1_value_payload_8[7:0]    ), //o
    .value_payload_9     (table_1_value_payload_9[7:0]    ), //o
    .value_payload_10    (table_1_value_payload_10[7:0]   ), //o
    .value_payload_11    (table_1_value_payload_11[7:0]   ), //o
    .value_payload_12    (table_1_value_payload_12[7:0]   ), //o
    .value_payload_13    (table_1_value_payload_13[7:0]   ), //o
    .value_payload_14    (table_1_value_payload_14[7:0]   ), //o
    .value_payload_15    (table_1_value_payload_15[7:0]   ), //o
    .clk                 (clk                             ), //i
    .reset               (reset                           )  //i
  );
  StreamDemux streamDemux_2 (
    .io_select                        (tmp_io_select_2[2:0]                              ), //i
    .io_input_valid                   (weightsAdapted_valid                              ), //i
    .io_input_ready                   (streamDemux_2_io_input_ready                      ), //o
    .io_input_payload_0_0_0_0         (weightsAdapted_payload_0_0_0_0[7:0]               ), //i
    .io_input_payload_0_0_0_1         (weightsAdapted_payload_0_0_0_1[7:0]               ), //i
    .io_input_payload_0_0_0_2         (weightsAdapted_payload_0_0_0_2[7:0]               ), //i
    .io_input_payload_0_0_0_3         (weightsAdapted_payload_0_0_0_3[7:0]               ), //i
    .io_input_payload_0_0_0_4         (weightsAdapted_payload_0_0_0_4[7:0]               ), //i
    .io_input_payload_0_0_0_5         (weightsAdapted_payload_0_0_0_5[7:0]               ), //i
    .io_input_payload_0_0_0_6         (weightsAdapted_payload_0_0_0_6[7:0]               ), //i
    .io_input_payload_0_0_0_7         (weightsAdapted_payload_0_0_0_7[7:0]               ), //i
    .io_input_payload_0_0_0_8         (weightsAdapted_payload_0_0_0_8[7:0]               ), //i
    .io_input_payload_0_0_0_9         (weightsAdapted_payload_0_0_0_9[7:0]               ), //i
    .io_input_payload_0_0_0_10        (weightsAdapted_payload_0_0_0_10[7:0]              ), //i
    .io_input_payload_0_0_0_11        (weightsAdapted_payload_0_0_0_11[7:0]              ), //i
    .io_input_payload_0_0_0_12        (weightsAdapted_payload_0_0_0_12[7:0]              ), //i
    .io_input_payload_0_0_0_13        (weightsAdapted_payload_0_0_0_13[7:0]              ), //i
    .io_input_payload_0_0_0_14        (weightsAdapted_payload_0_0_0_14[7:0]              ), //i
    .io_input_payload_0_0_0_15        (weightsAdapted_payload_0_0_0_15[7:0]              ), //i
    .io_input_payload_0_0_1_0         (weightsAdapted_payload_0_0_1_0[7:0]               ), //i
    .io_input_payload_0_0_1_1         (weightsAdapted_payload_0_0_1_1[7:0]               ), //i
    .io_input_payload_0_0_1_2         (weightsAdapted_payload_0_0_1_2[7:0]               ), //i
    .io_input_payload_0_0_1_3         (weightsAdapted_payload_0_0_1_3[7:0]               ), //i
    .io_input_payload_0_0_1_4         (weightsAdapted_payload_0_0_1_4[7:0]               ), //i
    .io_input_payload_0_0_1_5         (weightsAdapted_payload_0_0_1_5[7:0]               ), //i
    .io_input_payload_0_0_1_6         (weightsAdapted_payload_0_0_1_6[7:0]               ), //i
    .io_input_payload_0_0_1_7         (weightsAdapted_payload_0_0_1_7[7:0]               ), //i
    .io_input_payload_0_0_1_8         (weightsAdapted_payload_0_0_1_8[7:0]               ), //i
    .io_input_payload_0_0_1_9         (weightsAdapted_payload_0_0_1_9[7:0]               ), //i
    .io_input_payload_0_0_1_10        (weightsAdapted_payload_0_0_1_10[7:0]              ), //i
    .io_input_payload_0_0_1_11        (weightsAdapted_payload_0_0_1_11[7:0]              ), //i
    .io_input_payload_0_0_1_12        (weightsAdapted_payload_0_0_1_12[7:0]              ), //i
    .io_input_payload_0_0_1_13        (weightsAdapted_payload_0_0_1_13[7:0]              ), //i
    .io_input_payload_0_0_1_14        (weightsAdapted_payload_0_0_1_14[7:0]              ), //i
    .io_input_payload_0_0_1_15        (weightsAdapted_payload_0_0_1_15[7:0]              ), //i
    .io_input_payload_0_0_2_0         (weightsAdapted_payload_0_0_2_0[7:0]               ), //i
    .io_input_payload_0_0_2_1         (weightsAdapted_payload_0_0_2_1[7:0]               ), //i
    .io_input_payload_0_0_2_2         (weightsAdapted_payload_0_0_2_2[7:0]               ), //i
    .io_input_payload_0_0_2_3         (weightsAdapted_payload_0_0_2_3[7:0]               ), //i
    .io_input_payload_0_0_2_4         (weightsAdapted_payload_0_0_2_4[7:0]               ), //i
    .io_input_payload_0_0_2_5         (weightsAdapted_payload_0_0_2_5[7:0]               ), //i
    .io_input_payload_0_0_2_6         (weightsAdapted_payload_0_0_2_6[7:0]               ), //i
    .io_input_payload_0_0_2_7         (weightsAdapted_payload_0_0_2_7[7:0]               ), //i
    .io_input_payload_0_0_2_8         (weightsAdapted_payload_0_0_2_8[7:0]               ), //i
    .io_input_payload_0_0_2_9         (weightsAdapted_payload_0_0_2_9[7:0]               ), //i
    .io_input_payload_0_0_2_10        (weightsAdapted_payload_0_0_2_10[7:0]              ), //i
    .io_input_payload_0_0_2_11        (weightsAdapted_payload_0_0_2_11[7:0]              ), //i
    .io_input_payload_0_0_2_12        (weightsAdapted_payload_0_0_2_12[7:0]              ), //i
    .io_input_payload_0_0_2_13        (weightsAdapted_payload_0_0_2_13[7:0]              ), //i
    .io_input_payload_0_0_2_14        (weightsAdapted_payload_0_0_2_14[7:0]              ), //i
    .io_input_payload_0_0_2_15        (weightsAdapted_payload_0_0_2_15[7:0]              ), //i
    .io_input_payload_0_1_0_0         (weightsAdapted_payload_0_1_0_0[7:0]               ), //i
    .io_input_payload_0_1_0_1         (weightsAdapted_payload_0_1_0_1[7:0]               ), //i
    .io_input_payload_0_1_0_2         (weightsAdapted_payload_0_1_0_2[7:0]               ), //i
    .io_input_payload_0_1_0_3         (weightsAdapted_payload_0_1_0_3[7:0]               ), //i
    .io_input_payload_0_1_0_4         (weightsAdapted_payload_0_1_0_4[7:0]               ), //i
    .io_input_payload_0_1_0_5         (weightsAdapted_payload_0_1_0_5[7:0]               ), //i
    .io_input_payload_0_1_0_6         (weightsAdapted_payload_0_1_0_6[7:0]               ), //i
    .io_input_payload_0_1_0_7         (weightsAdapted_payload_0_1_0_7[7:0]               ), //i
    .io_input_payload_0_1_0_8         (weightsAdapted_payload_0_1_0_8[7:0]               ), //i
    .io_input_payload_0_1_0_9         (weightsAdapted_payload_0_1_0_9[7:0]               ), //i
    .io_input_payload_0_1_0_10        (weightsAdapted_payload_0_1_0_10[7:0]              ), //i
    .io_input_payload_0_1_0_11        (weightsAdapted_payload_0_1_0_11[7:0]              ), //i
    .io_input_payload_0_1_0_12        (weightsAdapted_payload_0_1_0_12[7:0]              ), //i
    .io_input_payload_0_1_0_13        (weightsAdapted_payload_0_1_0_13[7:0]              ), //i
    .io_input_payload_0_1_0_14        (weightsAdapted_payload_0_1_0_14[7:0]              ), //i
    .io_input_payload_0_1_0_15        (weightsAdapted_payload_0_1_0_15[7:0]              ), //i
    .io_input_payload_0_1_1_0         (weightsAdapted_payload_0_1_1_0[7:0]               ), //i
    .io_input_payload_0_1_1_1         (weightsAdapted_payload_0_1_1_1[7:0]               ), //i
    .io_input_payload_0_1_1_2         (weightsAdapted_payload_0_1_1_2[7:0]               ), //i
    .io_input_payload_0_1_1_3         (weightsAdapted_payload_0_1_1_3[7:0]               ), //i
    .io_input_payload_0_1_1_4         (weightsAdapted_payload_0_1_1_4[7:0]               ), //i
    .io_input_payload_0_1_1_5         (weightsAdapted_payload_0_1_1_5[7:0]               ), //i
    .io_input_payload_0_1_1_6         (weightsAdapted_payload_0_1_1_6[7:0]               ), //i
    .io_input_payload_0_1_1_7         (weightsAdapted_payload_0_1_1_7[7:0]               ), //i
    .io_input_payload_0_1_1_8         (weightsAdapted_payload_0_1_1_8[7:0]               ), //i
    .io_input_payload_0_1_1_9         (weightsAdapted_payload_0_1_1_9[7:0]               ), //i
    .io_input_payload_0_1_1_10        (weightsAdapted_payload_0_1_1_10[7:0]              ), //i
    .io_input_payload_0_1_1_11        (weightsAdapted_payload_0_1_1_11[7:0]              ), //i
    .io_input_payload_0_1_1_12        (weightsAdapted_payload_0_1_1_12[7:0]              ), //i
    .io_input_payload_0_1_1_13        (weightsAdapted_payload_0_1_1_13[7:0]              ), //i
    .io_input_payload_0_1_1_14        (weightsAdapted_payload_0_1_1_14[7:0]              ), //i
    .io_input_payload_0_1_1_15        (weightsAdapted_payload_0_1_1_15[7:0]              ), //i
    .io_input_payload_0_1_2_0         (weightsAdapted_payload_0_1_2_0[7:0]               ), //i
    .io_input_payload_0_1_2_1         (weightsAdapted_payload_0_1_2_1[7:0]               ), //i
    .io_input_payload_0_1_2_2         (weightsAdapted_payload_0_1_2_2[7:0]               ), //i
    .io_input_payload_0_1_2_3         (weightsAdapted_payload_0_1_2_3[7:0]               ), //i
    .io_input_payload_0_1_2_4         (weightsAdapted_payload_0_1_2_4[7:0]               ), //i
    .io_input_payload_0_1_2_5         (weightsAdapted_payload_0_1_2_5[7:0]               ), //i
    .io_input_payload_0_1_2_6         (weightsAdapted_payload_0_1_2_6[7:0]               ), //i
    .io_input_payload_0_1_2_7         (weightsAdapted_payload_0_1_2_7[7:0]               ), //i
    .io_input_payload_0_1_2_8         (weightsAdapted_payload_0_1_2_8[7:0]               ), //i
    .io_input_payload_0_1_2_9         (weightsAdapted_payload_0_1_2_9[7:0]               ), //i
    .io_input_payload_0_1_2_10        (weightsAdapted_payload_0_1_2_10[7:0]              ), //i
    .io_input_payload_0_1_2_11        (weightsAdapted_payload_0_1_2_11[7:0]              ), //i
    .io_input_payload_0_1_2_12        (weightsAdapted_payload_0_1_2_12[7:0]              ), //i
    .io_input_payload_0_1_2_13        (weightsAdapted_payload_0_1_2_13[7:0]              ), //i
    .io_input_payload_0_1_2_14        (weightsAdapted_payload_0_1_2_14[7:0]              ), //i
    .io_input_payload_0_1_2_15        (weightsAdapted_payload_0_1_2_15[7:0]              ), //i
    .io_input_payload_0_2_0_0         (weightsAdapted_payload_0_2_0_0[7:0]               ), //i
    .io_input_payload_0_2_0_1         (weightsAdapted_payload_0_2_0_1[7:0]               ), //i
    .io_input_payload_0_2_0_2         (weightsAdapted_payload_0_2_0_2[7:0]               ), //i
    .io_input_payload_0_2_0_3         (weightsAdapted_payload_0_2_0_3[7:0]               ), //i
    .io_input_payload_0_2_0_4         (weightsAdapted_payload_0_2_0_4[7:0]               ), //i
    .io_input_payload_0_2_0_5         (weightsAdapted_payload_0_2_0_5[7:0]               ), //i
    .io_input_payload_0_2_0_6         (weightsAdapted_payload_0_2_0_6[7:0]               ), //i
    .io_input_payload_0_2_0_7         (weightsAdapted_payload_0_2_0_7[7:0]               ), //i
    .io_input_payload_0_2_0_8         (weightsAdapted_payload_0_2_0_8[7:0]               ), //i
    .io_input_payload_0_2_0_9         (weightsAdapted_payload_0_2_0_9[7:0]               ), //i
    .io_input_payload_0_2_0_10        (weightsAdapted_payload_0_2_0_10[7:0]              ), //i
    .io_input_payload_0_2_0_11        (weightsAdapted_payload_0_2_0_11[7:0]              ), //i
    .io_input_payload_0_2_0_12        (weightsAdapted_payload_0_2_0_12[7:0]              ), //i
    .io_input_payload_0_2_0_13        (weightsAdapted_payload_0_2_0_13[7:0]              ), //i
    .io_input_payload_0_2_0_14        (weightsAdapted_payload_0_2_0_14[7:0]              ), //i
    .io_input_payload_0_2_0_15        (weightsAdapted_payload_0_2_0_15[7:0]              ), //i
    .io_input_payload_0_2_1_0         (weightsAdapted_payload_0_2_1_0[7:0]               ), //i
    .io_input_payload_0_2_1_1         (weightsAdapted_payload_0_2_1_1[7:0]               ), //i
    .io_input_payload_0_2_1_2         (weightsAdapted_payload_0_2_1_2[7:0]               ), //i
    .io_input_payload_0_2_1_3         (weightsAdapted_payload_0_2_1_3[7:0]               ), //i
    .io_input_payload_0_2_1_4         (weightsAdapted_payload_0_2_1_4[7:0]               ), //i
    .io_input_payload_0_2_1_5         (weightsAdapted_payload_0_2_1_5[7:0]               ), //i
    .io_input_payload_0_2_1_6         (weightsAdapted_payload_0_2_1_6[7:0]               ), //i
    .io_input_payload_0_2_1_7         (weightsAdapted_payload_0_2_1_7[7:0]               ), //i
    .io_input_payload_0_2_1_8         (weightsAdapted_payload_0_2_1_8[7:0]               ), //i
    .io_input_payload_0_2_1_9         (weightsAdapted_payload_0_2_1_9[7:0]               ), //i
    .io_input_payload_0_2_1_10        (weightsAdapted_payload_0_2_1_10[7:0]              ), //i
    .io_input_payload_0_2_1_11        (weightsAdapted_payload_0_2_1_11[7:0]              ), //i
    .io_input_payload_0_2_1_12        (weightsAdapted_payload_0_2_1_12[7:0]              ), //i
    .io_input_payload_0_2_1_13        (weightsAdapted_payload_0_2_1_13[7:0]              ), //i
    .io_input_payload_0_2_1_14        (weightsAdapted_payload_0_2_1_14[7:0]              ), //i
    .io_input_payload_0_2_1_15        (weightsAdapted_payload_0_2_1_15[7:0]              ), //i
    .io_input_payload_0_2_2_0         (weightsAdapted_payload_0_2_2_0[7:0]               ), //i
    .io_input_payload_0_2_2_1         (weightsAdapted_payload_0_2_2_1[7:0]               ), //i
    .io_input_payload_0_2_2_2         (weightsAdapted_payload_0_2_2_2[7:0]               ), //i
    .io_input_payload_0_2_2_3         (weightsAdapted_payload_0_2_2_3[7:0]               ), //i
    .io_input_payload_0_2_2_4         (weightsAdapted_payload_0_2_2_4[7:0]               ), //i
    .io_input_payload_0_2_2_5         (weightsAdapted_payload_0_2_2_5[7:0]               ), //i
    .io_input_payload_0_2_2_6         (weightsAdapted_payload_0_2_2_6[7:0]               ), //i
    .io_input_payload_0_2_2_7         (weightsAdapted_payload_0_2_2_7[7:0]               ), //i
    .io_input_payload_0_2_2_8         (weightsAdapted_payload_0_2_2_8[7:0]               ), //i
    .io_input_payload_0_2_2_9         (weightsAdapted_payload_0_2_2_9[7:0]               ), //i
    .io_input_payload_0_2_2_10        (weightsAdapted_payload_0_2_2_10[7:0]              ), //i
    .io_input_payload_0_2_2_11        (weightsAdapted_payload_0_2_2_11[7:0]              ), //i
    .io_input_payload_0_2_2_12        (weightsAdapted_payload_0_2_2_12[7:0]              ), //i
    .io_input_payload_0_2_2_13        (weightsAdapted_payload_0_2_2_13[7:0]              ), //i
    .io_input_payload_0_2_2_14        (weightsAdapted_payload_0_2_2_14[7:0]              ), //i
    .io_input_payload_0_2_2_15        (weightsAdapted_payload_0_2_2_15[7:0]              ), //i
    .io_input_payload_1_0_0_0         (weightsAdapted_payload_1_0_0_0[7:0]               ), //i
    .io_input_payload_1_0_0_1         (weightsAdapted_payload_1_0_0_1[7:0]               ), //i
    .io_input_payload_1_0_0_2         (weightsAdapted_payload_1_0_0_2[7:0]               ), //i
    .io_input_payload_1_0_0_3         (weightsAdapted_payload_1_0_0_3[7:0]               ), //i
    .io_input_payload_1_0_0_4         (weightsAdapted_payload_1_0_0_4[7:0]               ), //i
    .io_input_payload_1_0_0_5         (weightsAdapted_payload_1_0_0_5[7:0]               ), //i
    .io_input_payload_1_0_0_6         (weightsAdapted_payload_1_0_0_6[7:0]               ), //i
    .io_input_payload_1_0_0_7         (weightsAdapted_payload_1_0_0_7[7:0]               ), //i
    .io_input_payload_1_0_0_8         (weightsAdapted_payload_1_0_0_8[7:0]               ), //i
    .io_input_payload_1_0_0_9         (weightsAdapted_payload_1_0_0_9[7:0]               ), //i
    .io_input_payload_1_0_0_10        (weightsAdapted_payload_1_0_0_10[7:0]              ), //i
    .io_input_payload_1_0_0_11        (weightsAdapted_payload_1_0_0_11[7:0]              ), //i
    .io_input_payload_1_0_0_12        (weightsAdapted_payload_1_0_0_12[7:0]              ), //i
    .io_input_payload_1_0_0_13        (weightsAdapted_payload_1_0_0_13[7:0]              ), //i
    .io_input_payload_1_0_0_14        (weightsAdapted_payload_1_0_0_14[7:0]              ), //i
    .io_input_payload_1_0_0_15        (weightsAdapted_payload_1_0_0_15[7:0]              ), //i
    .io_input_payload_1_0_1_0         (weightsAdapted_payload_1_0_1_0[7:0]               ), //i
    .io_input_payload_1_0_1_1         (weightsAdapted_payload_1_0_1_1[7:0]               ), //i
    .io_input_payload_1_0_1_2         (weightsAdapted_payload_1_0_1_2[7:0]               ), //i
    .io_input_payload_1_0_1_3         (weightsAdapted_payload_1_0_1_3[7:0]               ), //i
    .io_input_payload_1_0_1_4         (weightsAdapted_payload_1_0_1_4[7:0]               ), //i
    .io_input_payload_1_0_1_5         (weightsAdapted_payload_1_0_1_5[7:0]               ), //i
    .io_input_payload_1_0_1_6         (weightsAdapted_payload_1_0_1_6[7:0]               ), //i
    .io_input_payload_1_0_1_7         (weightsAdapted_payload_1_0_1_7[7:0]               ), //i
    .io_input_payload_1_0_1_8         (weightsAdapted_payload_1_0_1_8[7:0]               ), //i
    .io_input_payload_1_0_1_9         (weightsAdapted_payload_1_0_1_9[7:0]               ), //i
    .io_input_payload_1_0_1_10        (weightsAdapted_payload_1_0_1_10[7:0]              ), //i
    .io_input_payload_1_0_1_11        (weightsAdapted_payload_1_0_1_11[7:0]              ), //i
    .io_input_payload_1_0_1_12        (weightsAdapted_payload_1_0_1_12[7:0]              ), //i
    .io_input_payload_1_0_1_13        (weightsAdapted_payload_1_0_1_13[7:0]              ), //i
    .io_input_payload_1_0_1_14        (weightsAdapted_payload_1_0_1_14[7:0]              ), //i
    .io_input_payload_1_0_1_15        (weightsAdapted_payload_1_0_1_15[7:0]              ), //i
    .io_input_payload_1_0_2_0         (weightsAdapted_payload_1_0_2_0[7:0]               ), //i
    .io_input_payload_1_0_2_1         (weightsAdapted_payload_1_0_2_1[7:0]               ), //i
    .io_input_payload_1_0_2_2         (weightsAdapted_payload_1_0_2_2[7:0]               ), //i
    .io_input_payload_1_0_2_3         (weightsAdapted_payload_1_0_2_3[7:0]               ), //i
    .io_input_payload_1_0_2_4         (weightsAdapted_payload_1_0_2_4[7:0]               ), //i
    .io_input_payload_1_0_2_5         (weightsAdapted_payload_1_0_2_5[7:0]               ), //i
    .io_input_payload_1_0_2_6         (weightsAdapted_payload_1_0_2_6[7:0]               ), //i
    .io_input_payload_1_0_2_7         (weightsAdapted_payload_1_0_2_7[7:0]               ), //i
    .io_input_payload_1_0_2_8         (weightsAdapted_payload_1_0_2_8[7:0]               ), //i
    .io_input_payload_1_0_2_9         (weightsAdapted_payload_1_0_2_9[7:0]               ), //i
    .io_input_payload_1_0_2_10        (weightsAdapted_payload_1_0_2_10[7:0]              ), //i
    .io_input_payload_1_0_2_11        (weightsAdapted_payload_1_0_2_11[7:0]              ), //i
    .io_input_payload_1_0_2_12        (weightsAdapted_payload_1_0_2_12[7:0]              ), //i
    .io_input_payload_1_0_2_13        (weightsAdapted_payload_1_0_2_13[7:0]              ), //i
    .io_input_payload_1_0_2_14        (weightsAdapted_payload_1_0_2_14[7:0]              ), //i
    .io_input_payload_1_0_2_15        (weightsAdapted_payload_1_0_2_15[7:0]              ), //i
    .io_input_payload_1_1_0_0         (weightsAdapted_payload_1_1_0_0[7:0]               ), //i
    .io_input_payload_1_1_0_1         (weightsAdapted_payload_1_1_0_1[7:0]               ), //i
    .io_input_payload_1_1_0_2         (weightsAdapted_payload_1_1_0_2[7:0]               ), //i
    .io_input_payload_1_1_0_3         (weightsAdapted_payload_1_1_0_3[7:0]               ), //i
    .io_input_payload_1_1_0_4         (weightsAdapted_payload_1_1_0_4[7:0]               ), //i
    .io_input_payload_1_1_0_5         (weightsAdapted_payload_1_1_0_5[7:0]               ), //i
    .io_input_payload_1_1_0_6         (weightsAdapted_payload_1_1_0_6[7:0]               ), //i
    .io_input_payload_1_1_0_7         (weightsAdapted_payload_1_1_0_7[7:0]               ), //i
    .io_input_payload_1_1_0_8         (weightsAdapted_payload_1_1_0_8[7:0]               ), //i
    .io_input_payload_1_1_0_9         (weightsAdapted_payload_1_1_0_9[7:0]               ), //i
    .io_input_payload_1_1_0_10        (weightsAdapted_payload_1_1_0_10[7:0]              ), //i
    .io_input_payload_1_1_0_11        (weightsAdapted_payload_1_1_0_11[7:0]              ), //i
    .io_input_payload_1_1_0_12        (weightsAdapted_payload_1_1_0_12[7:0]              ), //i
    .io_input_payload_1_1_0_13        (weightsAdapted_payload_1_1_0_13[7:0]              ), //i
    .io_input_payload_1_1_0_14        (weightsAdapted_payload_1_1_0_14[7:0]              ), //i
    .io_input_payload_1_1_0_15        (weightsAdapted_payload_1_1_0_15[7:0]              ), //i
    .io_input_payload_1_1_1_0         (weightsAdapted_payload_1_1_1_0[7:0]               ), //i
    .io_input_payload_1_1_1_1         (weightsAdapted_payload_1_1_1_1[7:0]               ), //i
    .io_input_payload_1_1_1_2         (weightsAdapted_payload_1_1_1_2[7:0]               ), //i
    .io_input_payload_1_1_1_3         (weightsAdapted_payload_1_1_1_3[7:0]               ), //i
    .io_input_payload_1_1_1_4         (weightsAdapted_payload_1_1_1_4[7:0]               ), //i
    .io_input_payload_1_1_1_5         (weightsAdapted_payload_1_1_1_5[7:0]               ), //i
    .io_input_payload_1_1_1_6         (weightsAdapted_payload_1_1_1_6[7:0]               ), //i
    .io_input_payload_1_1_1_7         (weightsAdapted_payload_1_1_1_7[7:0]               ), //i
    .io_input_payload_1_1_1_8         (weightsAdapted_payload_1_1_1_8[7:0]               ), //i
    .io_input_payload_1_1_1_9         (weightsAdapted_payload_1_1_1_9[7:0]               ), //i
    .io_input_payload_1_1_1_10        (weightsAdapted_payload_1_1_1_10[7:0]              ), //i
    .io_input_payload_1_1_1_11        (weightsAdapted_payload_1_1_1_11[7:0]              ), //i
    .io_input_payload_1_1_1_12        (weightsAdapted_payload_1_1_1_12[7:0]              ), //i
    .io_input_payload_1_1_1_13        (weightsAdapted_payload_1_1_1_13[7:0]              ), //i
    .io_input_payload_1_1_1_14        (weightsAdapted_payload_1_1_1_14[7:0]              ), //i
    .io_input_payload_1_1_1_15        (weightsAdapted_payload_1_1_1_15[7:0]              ), //i
    .io_input_payload_1_1_2_0         (weightsAdapted_payload_1_1_2_0[7:0]               ), //i
    .io_input_payload_1_1_2_1         (weightsAdapted_payload_1_1_2_1[7:0]               ), //i
    .io_input_payload_1_1_2_2         (weightsAdapted_payload_1_1_2_2[7:0]               ), //i
    .io_input_payload_1_1_2_3         (weightsAdapted_payload_1_1_2_3[7:0]               ), //i
    .io_input_payload_1_1_2_4         (weightsAdapted_payload_1_1_2_4[7:0]               ), //i
    .io_input_payload_1_1_2_5         (weightsAdapted_payload_1_1_2_5[7:0]               ), //i
    .io_input_payload_1_1_2_6         (weightsAdapted_payload_1_1_2_6[7:0]               ), //i
    .io_input_payload_1_1_2_7         (weightsAdapted_payload_1_1_2_7[7:0]               ), //i
    .io_input_payload_1_1_2_8         (weightsAdapted_payload_1_1_2_8[7:0]               ), //i
    .io_input_payload_1_1_2_9         (weightsAdapted_payload_1_1_2_9[7:0]               ), //i
    .io_input_payload_1_1_2_10        (weightsAdapted_payload_1_1_2_10[7:0]              ), //i
    .io_input_payload_1_1_2_11        (weightsAdapted_payload_1_1_2_11[7:0]              ), //i
    .io_input_payload_1_1_2_12        (weightsAdapted_payload_1_1_2_12[7:0]              ), //i
    .io_input_payload_1_1_2_13        (weightsAdapted_payload_1_1_2_13[7:0]              ), //i
    .io_input_payload_1_1_2_14        (weightsAdapted_payload_1_1_2_14[7:0]              ), //i
    .io_input_payload_1_1_2_15        (weightsAdapted_payload_1_1_2_15[7:0]              ), //i
    .io_input_payload_1_2_0_0         (weightsAdapted_payload_1_2_0_0[7:0]               ), //i
    .io_input_payload_1_2_0_1         (weightsAdapted_payload_1_2_0_1[7:0]               ), //i
    .io_input_payload_1_2_0_2         (weightsAdapted_payload_1_2_0_2[7:0]               ), //i
    .io_input_payload_1_2_0_3         (weightsAdapted_payload_1_2_0_3[7:0]               ), //i
    .io_input_payload_1_2_0_4         (weightsAdapted_payload_1_2_0_4[7:0]               ), //i
    .io_input_payload_1_2_0_5         (weightsAdapted_payload_1_2_0_5[7:0]               ), //i
    .io_input_payload_1_2_0_6         (weightsAdapted_payload_1_2_0_6[7:0]               ), //i
    .io_input_payload_1_2_0_7         (weightsAdapted_payload_1_2_0_7[7:0]               ), //i
    .io_input_payload_1_2_0_8         (weightsAdapted_payload_1_2_0_8[7:0]               ), //i
    .io_input_payload_1_2_0_9         (weightsAdapted_payload_1_2_0_9[7:0]               ), //i
    .io_input_payload_1_2_0_10        (weightsAdapted_payload_1_2_0_10[7:0]              ), //i
    .io_input_payload_1_2_0_11        (weightsAdapted_payload_1_2_0_11[7:0]              ), //i
    .io_input_payload_1_2_0_12        (weightsAdapted_payload_1_2_0_12[7:0]              ), //i
    .io_input_payload_1_2_0_13        (weightsAdapted_payload_1_2_0_13[7:0]              ), //i
    .io_input_payload_1_2_0_14        (weightsAdapted_payload_1_2_0_14[7:0]              ), //i
    .io_input_payload_1_2_0_15        (weightsAdapted_payload_1_2_0_15[7:0]              ), //i
    .io_input_payload_1_2_1_0         (weightsAdapted_payload_1_2_1_0[7:0]               ), //i
    .io_input_payload_1_2_1_1         (weightsAdapted_payload_1_2_1_1[7:0]               ), //i
    .io_input_payload_1_2_1_2         (weightsAdapted_payload_1_2_1_2[7:0]               ), //i
    .io_input_payload_1_2_1_3         (weightsAdapted_payload_1_2_1_3[7:0]               ), //i
    .io_input_payload_1_2_1_4         (weightsAdapted_payload_1_2_1_4[7:0]               ), //i
    .io_input_payload_1_2_1_5         (weightsAdapted_payload_1_2_1_5[7:0]               ), //i
    .io_input_payload_1_2_1_6         (weightsAdapted_payload_1_2_1_6[7:0]               ), //i
    .io_input_payload_1_2_1_7         (weightsAdapted_payload_1_2_1_7[7:0]               ), //i
    .io_input_payload_1_2_1_8         (weightsAdapted_payload_1_2_1_8[7:0]               ), //i
    .io_input_payload_1_2_1_9         (weightsAdapted_payload_1_2_1_9[7:0]               ), //i
    .io_input_payload_1_2_1_10        (weightsAdapted_payload_1_2_1_10[7:0]              ), //i
    .io_input_payload_1_2_1_11        (weightsAdapted_payload_1_2_1_11[7:0]              ), //i
    .io_input_payload_1_2_1_12        (weightsAdapted_payload_1_2_1_12[7:0]              ), //i
    .io_input_payload_1_2_1_13        (weightsAdapted_payload_1_2_1_13[7:0]              ), //i
    .io_input_payload_1_2_1_14        (weightsAdapted_payload_1_2_1_14[7:0]              ), //i
    .io_input_payload_1_2_1_15        (weightsAdapted_payload_1_2_1_15[7:0]              ), //i
    .io_input_payload_1_2_2_0         (weightsAdapted_payload_1_2_2_0[7:0]               ), //i
    .io_input_payload_1_2_2_1         (weightsAdapted_payload_1_2_2_1[7:0]               ), //i
    .io_input_payload_1_2_2_2         (weightsAdapted_payload_1_2_2_2[7:0]               ), //i
    .io_input_payload_1_2_2_3         (weightsAdapted_payload_1_2_2_3[7:0]               ), //i
    .io_input_payload_1_2_2_4         (weightsAdapted_payload_1_2_2_4[7:0]               ), //i
    .io_input_payload_1_2_2_5         (weightsAdapted_payload_1_2_2_5[7:0]               ), //i
    .io_input_payload_1_2_2_6         (weightsAdapted_payload_1_2_2_6[7:0]               ), //i
    .io_input_payload_1_2_2_7         (weightsAdapted_payload_1_2_2_7[7:0]               ), //i
    .io_input_payload_1_2_2_8         (weightsAdapted_payload_1_2_2_8[7:0]               ), //i
    .io_input_payload_1_2_2_9         (weightsAdapted_payload_1_2_2_9[7:0]               ), //i
    .io_input_payload_1_2_2_10        (weightsAdapted_payload_1_2_2_10[7:0]              ), //i
    .io_input_payload_1_2_2_11        (weightsAdapted_payload_1_2_2_11[7:0]              ), //i
    .io_input_payload_1_2_2_12        (weightsAdapted_payload_1_2_2_12[7:0]              ), //i
    .io_input_payload_1_2_2_13        (weightsAdapted_payload_1_2_2_13[7:0]              ), //i
    .io_input_payload_1_2_2_14        (weightsAdapted_payload_1_2_2_14[7:0]              ), //i
    .io_input_payload_1_2_2_15        (weightsAdapted_payload_1_2_2_15[7:0]              ), //i
    .io_outputs_0_valid               (streamDemux_2_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready               (weightFifo_0_push_ready                           ), //i
    .io_outputs_0_payload_0_0_0_0     (streamDemux_2_io_outputs_0_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_1     (streamDemux_2_io_outputs_0_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_2     (streamDemux_2_io_outputs_0_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_3     (streamDemux_2_io_outputs_0_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_4     (streamDemux_2_io_outputs_0_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_5     (streamDemux_2_io_outputs_0_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_6     (streamDemux_2_io_outputs_0_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_7     (streamDemux_2_io_outputs_0_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_8     (streamDemux_2_io_outputs_0_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_9     (streamDemux_2_io_outputs_0_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_0_payload_0_0_0_10    (streamDemux_2_io_outputs_0_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_0_payload_0_0_0_11    (streamDemux_2_io_outputs_0_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_0_payload_0_0_0_12    (streamDemux_2_io_outputs_0_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_0_payload_0_0_0_13    (streamDemux_2_io_outputs_0_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_0_payload_0_0_0_14    (streamDemux_2_io_outputs_0_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_0_payload_0_0_0_15    (streamDemux_2_io_outputs_0_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_0     (streamDemux_2_io_outputs_0_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_1     (streamDemux_2_io_outputs_0_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_2     (streamDemux_2_io_outputs_0_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_3     (streamDemux_2_io_outputs_0_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_4     (streamDemux_2_io_outputs_0_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_5     (streamDemux_2_io_outputs_0_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_6     (streamDemux_2_io_outputs_0_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_7     (streamDemux_2_io_outputs_0_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_8     (streamDemux_2_io_outputs_0_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_9     (streamDemux_2_io_outputs_0_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_0_payload_0_0_1_10    (streamDemux_2_io_outputs_0_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_11    (streamDemux_2_io_outputs_0_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_12    (streamDemux_2_io_outputs_0_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_13    (streamDemux_2_io_outputs_0_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_14    (streamDemux_2_io_outputs_0_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_0_payload_0_0_1_15    (streamDemux_2_io_outputs_0_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_0     (streamDemux_2_io_outputs_0_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_1     (streamDemux_2_io_outputs_0_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_2     (streamDemux_2_io_outputs_0_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_3     (streamDemux_2_io_outputs_0_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_4     (streamDemux_2_io_outputs_0_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_5     (streamDemux_2_io_outputs_0_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_6     (streamDemux_2_io_outputs_0_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_7     (streamDemux_2_io_outputs_0_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_8     (streamDemux_2_io_outputs_0_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_9     (streamDemux_2_io_outputs_0_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_0_payload_0_0_2_10    (streamDemux_2_io_outputs_0_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_11    (streamDemux_2_io_outputs_0_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_12    (streamDemux_2_io_outputs_0_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_13    (streamDemux_2_io_outputs_0_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_14    (streamDemux_2_io_outputs_0_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_0_payload_0_0_2_15    (streamDemux_2_io_outputs_0_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_0     (streamDemux_2_io_outputs_0_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_1     (streamDemux_2_io_outputs_0_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_2     (streamDemux_2_io_outputs_0_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_3     (streamDemux_2_io_outputs_0_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_4     (streamDemux_2_io_outputs_0_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_5     (streamDemux_2_io_outputs_0_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_6     (streamDemux_2_io_outputs_0_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_7     (streamDemux_2_io_outputs_0_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_8     (streamDemux_2_io_outputs_0_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_9     (streamDemux_2_io_outputs_0_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_0_payload_0_1_0_10    (streamDemux_2_io_outputs_0_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_11    (streamDemux_2_io_outputs_0_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_12    (streamDemux_2_io_outputs_0_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_13    (streamDemux_2_io_outputs_0_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_14    (streamDemux_2_io_outputs_0_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_0_payload_0_1_0_15    (streamDemux_2_io_outputs_0_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_0     (streamDemux_2_io_outputs_0_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_1     (streamDemux_2_io_outputs_0_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_2     (streamDemux_2_io_outputs_0_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_3     (streamDemux_2_io_outputs_0_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_4     (streamDemux_2_io_outputs_0_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_5     (streamDemux_2_io_outputs_0_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_6     (streamDemux_2_io_outputs_0_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_7     (streamDemux_2_io_outputs_0_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_8     (streamDemux_2_io_outputs_0_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_9     (streamDemux_2_io_outputs_0_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_0_payload_0_1_1_10    (streamDemux_2_io_outputs_0_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_11    (streamDemux_2_io_outputs_0_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_12    (streamDemux_2_io_outputs_0_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_13    (streamDemux_2_io_outputs_0_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_14    (streamDemux_2_io_outputs_0_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_0_payload_0_1_1_15    (streamDemux_2_io_outputs_0_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_0     (streamDemux_2_io_outputs_0_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_1     (streamDemux_2_io_outputs_0_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_2     (streamDemux_2_io_outputs_0_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_3     (streamDemux_2_io_outputs_0_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_4     (streamDemux_2_io_outputs_0_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_5     (streamDemux_2_io_outputs_0_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_6     (streamDemux_2_io_outputs_0_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_7     (streamDemux_2_io_outputs_0_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_8     (streamDemux_2_io_outputs_0_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_9     (streamDemux_2_io_outputs_0_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_0_payload_0_1_2_10    (streamDemux_2_io_outputs_0_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_11    (streamDemux_2_io_outputs_0_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_12    (streamDemux_2_io_outputs_0_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_13    (streamDemux_2_io_outputs_0_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_14    (streamDemux_2_io_outputs_0_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_0_payload_0_1_2_15    (streamDemux_2_io_outputs_0_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_0     (streamDemux_2_io_outputs_0_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_1     (streamDemux_2_io_outputs_0_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_2     (streamDemux_2_io_outputs_0_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_3     (streamDemux_2_io_outputs_0_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_4     (streamDemux_2_io_outputs_0_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_5     (streamDemux_2_io_outputs_0_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_6     (streamDemux_2_io_outputs_0_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_7     (streamDemux_2_io_outputs_0_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_8     (streamDemux_2_io_outputs_0_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_9     (streamDemux_2_io_outputs_0_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_0_payload_0_2_0_10    (streamDemux_2_io_outputs_0_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_11    (streamDemux_2_io_outputs_0_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_12    (streamDemux_2_io_outputs_0_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_13    (streamDemux_2_io_outputs_0_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_14    (streamDemux_2_io_outputs_0_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_0_payload_0_2_0_15    (streamDemux_2_io_outputs_0_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_0     (streamDemux_2_io_outputs_0_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_1     (streamDemux_2_io_outputs_0_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_2     (streamDemux_2_io_outputs_0_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_3     (streamDemux_2_io_outputs_0_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_4     (streamDemux_2_io_outputs_0_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_5     (streamDemux_2_io_outputs_0_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_6     (streamDemux_2_io_outputs_0_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_7     (streamDemux_2_io_outputs_0_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_8     (streamDemux_2_io_outputs_0_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_9     (streamDemux_2_io_outputs_0_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_0_payload_0_2_1_10    (streamDemux_2_io_outputs_0_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_11    (streamDemux_2_io_outputs_0_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_12    (streamDemux_2_io_outputs_0_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_13    (streamDemux_2_io_outputs_0_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_14    (streamDemux_2_io_outputs_0_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_0_payload_0_2_1_15    (streamDemux_2_io_outputs_0_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_0     (streamDemux_2_io_outputs_0_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_1     (streamDemux_2_io_outputs_0_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_2     (streamDemux_2_io_outputs_0_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_3     (streamDemux_2_io_outputs_0_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_4     (streamDemux_2_io_outputs_0_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_5     (streamDemux_2_io_outputs_0_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_6     (streamDemux_2_io_outputs_0_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_7     (streamDemux_2_io_outputs_0_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_8     (streamDemux_2_io_outputs_0_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_9     (streamDemux_2_io_outputs_0_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_0_payload_0_2_2_10    (streamDemux_2_io_outputs_0_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_11    (streamDemux_2_io_outputs_0_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_12    (streamDemux_2_io_outputs_0_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_13    (streamDemux_2_io_outputs_0_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_14    (streamDemux_2_io_outputs_0_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_0_payload_0_2_2_15    (streamDemux_2_io_outputs_0_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_0     (streamDemux_2_io_outputs_0_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_1     (streamDemux_2_io_outputs_0_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_2     (streamDemux_2_io_outputs_0_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_3     (streamDemux_2_io_outputs_0_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_4     (streamDemux_2_io_outputs_0_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_5     (streamDemux_2_io_outputs_0_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_6     (streamDemux_2_io_outputs_0_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_7     (streamDemux_2_io_outputs_0_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_8     (streamDemux_2_io_outputs_0_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_9     (streamDemux_2_io_outputs_0_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_0_payload_1_0_0_10    (streamDemux_2_io_outputs_0_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_11    (streamDemux_2_io_outputs_0_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_12    (streamDemux_2_io_outputs_0_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_13    (streamDemux_2_io_outputs_0_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_14    (streamDemux_2_io_outputs_0_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_0_payload_1_0_0_15    (streamDemux_2_io_outputs_0_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_0     (streamDemux_2_io_outputs_0_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_1     (streamDemux_2_io_outputs_0_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_2     (streamDemux_2_io_outputs_0_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_3     (streamDemux_2_io_outputs_0_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_4     (streamDemux_2_io_outputs_0_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_5     (streamDemux_2_io_outputs_0_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_6     (streamDemux_2_io_outputs_0_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_7     (streamDemux_2_io_outputs_0_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_8     (streamDemux_2_io_outputs_0_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_9     (streamDemux_2_io_outputs_0_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_0_payload_1_0_1_10    (streamDemux_2_io_outputs_0_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_11    (streamDemux_2_io_outputs_0_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_12    (streamDemux_2_io_outputs_0_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_13    (streamDemux_2_io_outputs_0_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_14    (streamDemux_2_io_outputs_0_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_0_payload_1_0_1_15    (streamDemux_2_io_outputs_0_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_0     (streamDemux_2_io_outputs_0_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_1     (streamDemux_2_io_outputs_0_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_2     (streamDemux_2_io_outputs_0_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_3     (streamDemux_2_io_outputs_0_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_4     (streamDemux_2_io_outputs_0_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_5     (streamDemux_2_io_outputs_0_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_6     (streamDemux_2_io_outputs_0_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_7     (streamDemux_2_io_outputs_0_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_8     (streamDemux_2_io_outputs_0_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_9     (streamDemux_2_io_outputs_0_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_0_payload_1_0_2_10    (streamDemux_2_io_outputs_0_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_11    (streamDemux_2_io_outputs_0_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_12    (streamDemux_2_io_outputs_0_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_13    (streamDemux_2_io_outputs_0_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_14    (streamDemux_2_io_outputs_0_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_0_payload_1_0_2_15    (streamDemux_2_io_outputs_0_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_0     (streamDemux_2_io_outputs_0_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_1     (streamDemux_2_io_outputs_0_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_2     (streamDemux_2_io_outputs_0_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_3     (streamDemux_2_io_outputs_0_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_4     (streamDemux_2_io_outputs_0_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_5     (streamDemux_2_io_outputs_0_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_6     (streamDemux_2_io_outputs_0_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_7     (streamDemux_2_io_outputs_0_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_8     (streamDemux_2_io_outputs_0_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_9     (streamDemux_2_io_outputs_0_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_0_payload_1_1_0_10    (streamDemux_2_io_outputs_0_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_11    (streamDemux_2_io_outputs_0_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_12    (streamDemux_2_io_outputs_0_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_13    (streamDemux_2_io_outputs_0_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_14    (streamDemux_2_io_outputs_0_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_0_payload_1_1_0_15    (streamDemux_2_io_outputs_0_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_0     (streamDemux_2_io_outputs_0_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_1     (streamDemux_2_io_outputs_0_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_2     (streamDemux_2_io_outputs_0_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_3     (streamDemux_2_io_outputs_0_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_4     (streamDemux_2_io_outputs_0_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_5     (streamDemux_2_io_outputs_0_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_6     (streamDemux_2_io_outputs_0_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_7     (streamDemux_2_io_outputs_0_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_8     (streamDemux_2_io_outputs_0_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_9     (streamDemux_2_io_outputs_0_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_0_payload_1_1_1_10    (streamDemux_2_io_outputs_0_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_11    (streamDemux_2_io_outputs_0_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_12    (streamDemux_2_io_outputs_0_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_13    (streamDemux_2_io_outputs_0_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_14    (streamDemux_2_io_outputs_0_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_0_payload_1_1_1_15    (streamDemux_2_io_outputs_0_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_0     (streamDemux_2_io_outputs_0_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_1     (streamDemux_2_io_outputs_0_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_2     (streamDemux_2_io_outputs_0_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_3     (streamDemux_2_io_outputs_0_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_4     (streamDemux_2_io_outputs_0_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_5     (streamDemux_2_io_outputs_0_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_6     (streamDemux_2_io_outputs_0_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_7     (streamDemux_2_io_outputs_0_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_8     (streamDemux_2_io_outputs_0_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_9     (streamDemux_2_io_outputs_0_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_0_payload_1_1_2_10    (streamDemux_2_io_outputs_0_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_11    (streamDemux_2_io_outputs_0_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_12    (streamDemux_2_io_outputs_0_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_13    (streamDemux_2_io_outputs_0_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_14    (streamDemux_2_io_outputs_0_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_0_payload_1_1_2_15    (streamDemux_2_io_outputs_0_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_0     (streamDemux_2_io_outputs_0_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_1     (streamDemux_2_io_outputs_0_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_2     (streamDemux_2_io_outputs_0_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_3     (streamDemux_2_io_outputs_0_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_4     (streamDemux_2_io_outputs_0_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_5     (streamDemux_2_io_outputs_0_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_6     (streamDemux_2_io_outputs_0_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_7     (streamDemux_2_io_outputs_0_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_8     (streamDemux_2_io_outputs_0_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_9     (streamDemux_2_io_outputs_0_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_0_payload_1_2_0_10    (streamDemux_2_io_outputs_0_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_11    (streamDemux_2_io_outputs_0_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_12    (streamDemux_2_io_outputs_0_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_13    (streamDemux_2_io_outputs_0_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_14    (streamDemux_2_io_outputs_0_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_0_payload_1_2_0_15    (streamDemux_2_io_outputs_0_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_0     (streamDemux_2_io_outputs_0_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_1     (streamDemux_2_io_outputs_0_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_2     (streamDemux_2_io_outputs_0_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_3     (streamDemux_2_io_outputs_0_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_4     (streamDemux_2_io_outputs_0_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_5     (streamDemux_2_io_outputs_0_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_6     (streamDemux_2_io_outputs_0_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_7     (streamDemux_2_io_outputs_0_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_8     (streamDemux_2_io_outputs_0_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_9     (streamDemux_2_io_outputs_0_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_0_payload_1_2_1_10    (streamDemux_2_io_outputs_0_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_11    (streamDemux_2_io_outputs_0_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_12    (streamDemux_2_io_outputs_0_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_13    (streamDemux_2_io_outputs_0_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_14    (streamDemux_2_io_outputs_0_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_0_payload_1_2_1_15    (streamDemux_2_io_outputs_0_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_0     (streamDemux_2_io_outputs_0_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_1     (streamDemux_2_io_outputs_0_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_2     (streamDemux_2_io_outputs_0_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_3     (streamDemux_2_io_outputs_0_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_4     (streamDemux_2_io_outputs_0_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_5     (streamDemux_2_io_outputs_0_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_6     (streamDemux_2_io_outputs_0_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_7     (streamDemux_2_io_outputs_0_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_8     (streamDemux_2_io_outputs_0_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_9     (streamDemux_2_io_outputs_0_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_0_payload_1_2_2_10    (streamDemux_2_io_outputs_0_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_11    (streamDemux_2_io_outputs_0_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_12    (streamDemux_2_io_outputs_0_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_13    (streamDemux_2_io_outputs_0_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_14    (streamDemux_2_io_outputs_0_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_0_payload_1_2_2_15    (streamDemux_2_io_outputs_0_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_1_valid               (streamDemux_2_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready               (weightFifo_1_push_ready                           ), //i
    .io_outputs_1_payload_0_0_0_0     (streamDemux_2_io_outputs_1_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_1     (streamDemux_2_io_outputs_1_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_2     (streamDemux_2_io_outputs_1_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_3     (streamDemux_2_io_outputs_1_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_4     (streamDemux_2_io_outputs_1_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_5     (streamDemux_2_io_outputs_1_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_6     (streamDemux_2_io_outputs_1_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_7     (streamDemux_2_io_outputs_1_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_8     (streamDemux_2_io_outputs_1_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_9     (streamDemux_2_io_outputs_1_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_1_payload_0_0_0_10    (streamDemux_2_io_outputs_1_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_1_payload_0_0_0_11    (streamDemux_2_io_outputs_1_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_1_payload_0_0_0_12    (streamDemux_2_io_outputs_1_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_1_payload_0_0_0_13    (streamDemux_2_io_outputs_1_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_1_payload_0_0_0_14    (streamDemux_2_io_outputs_1_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_1_payload_0_0_0_15    (streamDemux_2_io_outputs_1_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_0     (streamDemux_2_io_outputs_1_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_1     (streamDemux_2_io_outputs_1_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_2     (streamDemux_2_io_outputs_1_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_3     (streamDemux_2_io_outputs_1_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_4     (streamDemux_2_io_outputs_1_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_5     (streamDemux_2_io_outputs_1_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_6     (streamDemux_2_io_outputs_1_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_7     (streamDemux_2_io_outputs_1_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_8     (streamDemux_2_io_outputs_1_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_9     (streamDemux_2_io_outputs_1_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_1_payload_0_0_1_10    (streamDemux_2_io_outputs_1_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_11    (streamDemux_2_io_outputs_1_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_12    (streamDemux_2_io_outputs_1_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_13    (streamDemux_2_io_outputs_1_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_14    (streamDemux_2_io_outputs_1_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_1_payload_0_0_1_15    (streamDemux_2_io_outputs_1_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_0     (streamDemux_2_io_outputs_1_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_1     (streamDemux_2_io_outputs_1_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_2     (streamDemux_2_io_outputs_1_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_3     (streamDemux_2_io_outputs_1_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_4     (streamDemux_2_io_outputs_1_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_5     (streamDemux_2_io_outputs_1_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_6     (streamDemux_2_io_outputs_1_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_7     (streamDemux_2_io_outputs_1_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_8     (streamDemux_2_io_outputs_1_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_9     (streamDemux_2_io_outputs_1_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_1_payload_0_0_2_10    (streamDemux_2_io_outputs_1_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_11    (streamDemux_2_io_outputs_1_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_12    (streamDemux_2_io_outputs_1_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_13    (streamDemux_2_io_outputs_1_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_14    (streamDemux_2_io_outputs_1_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_1_payload_0_0_2_15    (streamDemux_2_io_outputs_1_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_0     (streamDemux_2_io_outputs_1_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_1     (streamDemux_2_io_outputs_1_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_2     (streamDemux_2_io_outputs_1_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_3     (streamDemux_2_io_outputs_1_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_4     (streamDemux_2_io_outputs_1_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_5     (streamDemux_2_io_outputs_1_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_6     (streamDemux_2_io_outputs_1_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_7     (streamDemux_2_io_outputs_1_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_8     (streamDemux_2_io_outputs_1_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_9     (streamDemux_2_io_outputs_1_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_1_payload_0_1_0_10    (streamDemux_2_io_outputs_1_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_11    (streamDemux_2_io_outputs_1_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_12    (streamDemux_2_io_outputs_1_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_13    (streamDemux_2_io_outputs_1_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_14    (streamDemux_2_io_outputs_1_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_1_payload_0_1_0_15    (streamDemux_2_io_outputs_1_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_0     (streamDemux_2_io_outputs_1_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_1     (streamDemux_2_io_outputs_1_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_2     (streamDemux_2_io_outputs_1_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_3     (streamDemux_2_io_outputs_1_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_4     (streamDemux_2_io_outputs_1_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_5     (streamDemux_2_io_outputs_1_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_6     (streamDemux_2_io_outputs_1_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_7     (streamDemux_2_io_outputs_1_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_8     (streamDemux_2_io_outputs_1_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_9     (streamDemux_2_io_outputs_1_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_1_payload_0_1_1_10    (streamDemux_2_io_outputs_1_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_11    (streamDemux_2_io_outputs_1_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_12    (streamDemux_2_io_outputs_1_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_13    (streamDemux_2_io_outputs_1_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_14    (streamDemux_2_io_outputs_1_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_1_payload_0_1_1_15    (streamDemux_2_io_outputs_1_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_0     (streamDemux_2_io_outputs_1_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_1     (streamDemux_2_io_outputs_1_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_2     (streamDemux_2_io_outputs_1_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_3     (streamDemux_2_io_outputs_1_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_4     (streamDemux_2_io_outputs_1_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_5     (streamDemux_2_io_outputs_1_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_6     (streamDemux_2_io_outputs_1_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_7     (streamDemux_2_io_outputs_1_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_8     (streamDemux_2_io_outputs_1_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_9     (streamDemux_2_io_outputs_1_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_1_payload_0_1_2_10    (streamDemux_2_io_outputs_1_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_11    (streamDemux_2_io_outputs_1_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_12    (streamDemux_2_io_outputs_1_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_13    (streamDemux_2_io_outputs_1_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_14    (streamDemux_2_io_outputs_1_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_1_payload_0_1_2_15    (streamDemux_2_io_outputs_1_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_0     (streamDemux_2_io_outputs_1_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_1     (streamDemux_2_io_outputs_1_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_2     (streamDemux_2_io_outputs_1_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_3     (streamDemux_2_io_outputs_1_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_4     (streamDemux_2_io_outputs_1_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_5     (streamDemux_2_io_outputs_1_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_6     (streamDemux_2_io_outputs_1_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_7     (streamDemux_2_io_outputs_1_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_8     (streamDemux_2_io_outputs_1_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_9     (streamDemux_2_io_outputs_1_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_1_payload_0_2_0_10    (streamDemux_2_io_outputs_1_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_11    (streamDemux_2_io_outputs_1_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_12    (streamDemux_2_io_outputs_1_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_13    (streamDemux_2_io_outputs_1_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_14    (streamDemux_2_io_outputs_1_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_1_payload_0_2_0_15    (streamDemux_2_io_outputs_1_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_0     (streamDemux_2_io_outputs_1_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_1     (streamDemux_2_io_outputs_1_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_2     (streamDemux_2_io_outputs_1_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_3     (streamDemux_2_io_outputs_1_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_4     (streamDemux_2_io_outputs_1_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_5     (streamDemux_2_io_outputs_1_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_6     (streamDemux_2_io_outputs_1_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_7     (streamDemux_2_io_outputs_1_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_8     (streamDemux_2_io_outputs_1_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_9     (streamDemux_2_io_outputs_1_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_1_payload_0_2_1_10    (streamDemux_2_io_outputs_1_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_11    (streamDemux_2_io_outputs_1_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_12    (streamDemux_2_io_outputs_1_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_13    (streamDemux_2_io_outputs_1_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_14    (streamDemux_2_io_outputs_1_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_1_payload_0_2_1_15    (streamDemux_2_io_outputs_1_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_0     (streamDemux_2_io_outputs_1_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_1     (streamDemux_2_io_outputs_1_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_2     (streamDemux_2_io_outputs_1_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_3     (streamDemux_2_io_outputs_1_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_4     (streamDemux_2_io_outputs_1_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_5     (streamDemux_2_io_outputs_1_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_6     (streamDemux_2_io_outputs_1_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_7     (streamDemux_2_io_outputs_1_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_8     (streamDemux_2_io_outputs_1_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_9     (streamDemux_2_io_outputs_1_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_1_payload_0_2_2_10    (streamDemux_2_io_outputs_1_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_11    (streamDemux_2_io_outputs_1_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_12    (streamDemux_2_io_outputs_1_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_13    (streamDemux_2_io_outputs_1_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_14    (streamDemux_2_io_outputs_1_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_1_payload_0_2_2_15    (streamDemux_2_io_outputs_1_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_0     (streamDemux_2_io_outputs_1_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_1     (streamDemux_2_io_outputs_1_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_2     (streamDemux_2_io_outputs_1_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_3     (streamDemux_2_io_outputs_1_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_4     (streamDemux_2_io_outputs_1_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_5     (streamDemux_2_io_outputs_1_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_6     (streamDemux_2_io_outputs_1_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_7     (streamDemux_2_io_outputs_1_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_8     (streamDemux_2_io_outputs_1_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_9     (streamDemux_2_io_outputs_1_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_1_payload_1_0_0_10    (streamDemux_2_io_outputs_1_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_11    (streamDemux_2_io_outputs_1_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_12    (streamDemux_2_io_outputs_1_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_13    (streamDemux_2_io_outputs_1_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_14    (streamDemux_2_io_outputs_1_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_1_payload_1_0_0_15    (streamDemux_2_io_outputs_1_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_0     (streamDemux_2_io_outputs_1_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_1     (streamDemux_2_io_outputs_1_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_2     (streamDemux_2_io_outputs_1_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_3     (streamDemux_2_io_outputs_1_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_4     (streamDemux_2_io_outputs_1_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_5     (streamDemux_2_io_outputs_1_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_6     (streamDemux_2_io_outputs_1_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_7     (streamDemux_2_io_outputs_1_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_8     (streamDemux_2_io_outputs_1_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_9     (streamDemux_2_io_outputs_1_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_1_payload_1_0_1_10    (streamDemux_2_io_outputs_1_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_11    (streamDemux_2_io_outputs_1_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_12    (streamDemux_2_io_outputs_1_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_13    (streamDemux_2_io_outputs_1_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_14    (streamDemux_2_io_outputs_1_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_1_payload_1_0_1_15    (streamDemux_2_io_outputs_1_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_0     (streamDemux_2_io_outputs_1_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_1     (streamDemux_2_io_outputs_1_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_2     (streamDemux_2_io_outputs_1_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_3     (streamDemux_2_io_outputs_1_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_4     (streamDemux_2_io_outputs_1_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_5     (streamDemux_2_io_outputs_1_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_6     (streamDemux_2_io_outputs_1_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_7     (streamDemux_2_io_outputs_1_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_8     (streamDemux_2_io_outputs_1_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_9     (streamDemux_2_io_outputs_1_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_1_payload_1_0_2_10    (streamDemux_2_io_outputs_1_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_11    (streamDemux_2_io_outputs_1_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_12    (streamDemux_2_io_outputs_1_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_13    (streamDemux_2_io_outputs_1_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_14    (streamDemux_2_io_outputs_1_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_1_payload_1_0_2_15    (streamDemux_2_io_outputs_1_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_0     (streamDemux_2_io_outputs_1_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_1     (streamDemux_2_io_outputs_1_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_2     (streamDemux_2_io_outputs_1_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_3     (streamDemux_2_io_outputs_1_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_4     (streamDemux_2_io_outputs_1_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_5     (streamDemux_2_io_outputs_1_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_6     (streamDemux_2_io_outputs_1_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_7     (streamDemux_2_io_outputs_1_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_8     (streamDemux_2_io_outputs_1_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_9     (streamDemux_2_io_outputs_1_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_1_payload_1_1_0_10    (streamDemux_2_io_outputs_1_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_11    (streamDemux_2_io_outputs_1_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_12    (streamDemux_2_io_outputs_1_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_13    (streamDemux_2_io_outputs_1_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_14    (streamDemux_2_io_outputs_1_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_1_payload_1_1_0_15    (streamDemux_2_io_outputs_1_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_0     (streamDemux_2_io_outputs_1_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_1     (streamDemux_2_io_outputs_1_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_2     (streamDemux_2_io_outputs_1_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_3     (streamDemux_2_io_outputs_1_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_4     (streamDemux_2_io_outputs_1_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_5     (streamDemux_2_io_outputs_1_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_6     (streamDemux_2_io_outputs_1_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_7     (streamDemux_2_io_outputs_1_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_8     (streamDemux_2_io_outputs_1_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_9     (streamDemux_2_io_outputs_1_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_1_payload_1_1_1_10    (streamDemux_2_io_outputs_1_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_11    (streamDemux_2_io_outputs_1_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_12    (streamDemux_2_io_outputs_1_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_13    (streamDemux_2_io_outputs_1_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_14    (streamDemux_2_io_outputs_1_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_1_payload_1_1_1_15    (streamDemux_2_io_outputs_1_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_0     (streamDemux_2_io_outputs_1_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_1     (streamDemux_2_io_outputs_1_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_2     (streamDemux_2_io_outputs_1_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_3     (streamDemux_2_io_outputs_1_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_4     (streamDemux_2_io_outputs_1_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_5     (streamDemux_2_io_outputs_1_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_6     (streamDemux_2_io_outputs_1_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_7     (streamDemux_2_io_outputs_1_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_8     (streamDemux_2_io_outputs_1_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_9     (streamDemux_2_io_outputs_1_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_1_payload_1_1_2_10    (streamDemux_2_io_outputs_1_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_11    (streamDemux_2_io_outputs_1_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_12    (streamDemux_2_io_outputs_1_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_13    (streamDemux_2_io_outputs_1_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_14    (streamDemux_2_io_outputs_1_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_1_payload_1_1_2_15    (streamDemux_2_io_outputs_1_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_0     (streamDemux_2_io_outputs_1_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_1     (streamDemux_2_io_outputs_1_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_2     (streamDemux_2_io_outputs_1_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_3     (streamDemux_2_io_outputs_1_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_4     (streamDemux_2_io_outputs_1_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_5     (streamDemux_2_io_outputs_1_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_6     (streamDemux_2_io_outputs_1_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_7     (streamDemux_2_io_outputs_1_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_8     (streamDemux_2_io_outputs_1_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_9     (streamDemux_2_io_outputs_1_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_1_payload_1_2_0_10    (streamDemux_2_io_outputs_1_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_11    (streamDemux_2_io_outputs_1_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_12    (streamDemux_2_io_outputs_1_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_13    (streamDemux_2_io_outputs_1_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_14    (streamDemux_2_io_outputs_1_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_1_payload_1_2_0_15    (streamDemux_2_io_outputs_1_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_0     (streamDemux_2_io_outputs_1_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_1     (streamDemux_2_io_outputs_1_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_2     (streamDemux_2_io_outputs_1_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_3     (streamDemux_2_io_outputs_1_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_4     (streamDemux_2_io_outputs_1_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_5     (streamDemux_2_io_outputs_1_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_6     (streamDemux_2_io_outputs_1_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_7     (streamDemux_2_io_outputs_1_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_8     (streamDemux_2_io_outputs_1_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_9     (streamDemux_2_io_outputs_1_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_1_payload_1_2_1_10    (streamDemux_2_io_outputs_1_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_11    (streamDemux_2_io_outputs_1_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_12    (streamDemux_2_io_outputs_1_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_13    (streamDemux_2_io_outputs_1_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_14    (streamDemux_2_io_outputs_1_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_1_payload_1_2_1_15    (streamDemux_2_io_outputs_1_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_0     (streamDemux_2_io_outputs_1_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_1     (streamDemux_2_io_outputs_1_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_2     (streamDemux_2_io_outputs_1_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_3     (streamDemux_2_io_outputs_1_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_4     (streamDemux_2_io_outputs_1_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_5     (streamDemux_2_io_outputs_1_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_6     (streamDemux_2_io_outputs_1_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_7     (streamDemux_2_io_outputs_1_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_8     (streamDemux_2_io_outputs_1_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_9     (streamDemux_2_io_outputs_1_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_1_payload_1_2_2_10    (streamDemux_2_io_outputs_1_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_11    (streamDemux_2_io_outputs_1_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_12    (streamDemux_2_io_outputs_1_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_13    (streamDemux_2_io_outputs_1_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_14    (streamDemux_2_io_outputs_1_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_1_payload_1_2_2_15    (streamDemux_2_io_outputs_1_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_2_valid               (streamDemux_2_io_outputs_2_valid                  ), //o
    .io_outputs_2_ready               (weightFifo_2_push_ready                           ), //i
    .io_outputs_2_payload_0_0_0_0     (streamDemux_2_io_outputs_2_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_1     (streamDemux_2_io_outputs_2_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_2     (streamDemux_2_io_outputs_2_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_3     (streamDemux_2_io_outputs_2_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_4     (streamDemux_2_io_outputs_2_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_5     (streamDemux_2_io_outputs_2_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_6     (streamDemux_2_io_outputs_2_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_7     (streamDemux_2_io_outputs_2_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_8     (streamDemux_2_io_outputs_2_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_9     (streamDemux_2_io_outputs_2_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_2_payload_0_0_0_10    (streamDemux_2_io_outputs_2_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_2_payload_0_0_0_11    (streamDemux_2_io_outputs_2_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_2_payload_0_0_0_12    (streamDemux_2_io_outputs_2_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_2_payload_0_0_0_13    (streamDemux_2_io_outputs_2_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_2_payload_0_0_0_14    (streamDemux_2_io_outputs_2_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_2_payload_0_0_0_15    (streamDemux_2_io_outputs_2_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_0     (streamDemux_2_io_outputs_2_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_1     (streamDemux_2_io_outputs_2_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_2     (streamDemux_2_io_outputs_2_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_3     (streamDemux_2_io_outputs_2_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_4     (streamDemux_2_io_outputs_2_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_5     (streamDemux_2_io_outputs_2_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_6     (streamDemux_2_io_outputs_2_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_7     (streamDemux_2_io_outputs_2_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_8     (streamDemux_2_io_outputs_2_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_9     (streamDemux_2_io_outputs_2_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_2_payload_0_0_1_10    (streamDemux_2_io_outputs_2_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_11    (streamDemux_2_io_outputs_2_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_12    (streamDemux_2_io_outputs_2_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_13    (streamDemux_2_io_outputs_2_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_14    (streamDemux_2_io_outputs_2_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_2_payload_0_0_1_15    (streamDemux_2_io_outputs_2_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_0     (streamDemux_2_io_outputs_2_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_1     (streamDemux_2_io_outputs_2_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_2     (streamDemux_2_io_outputs_2_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_3     (streamDemux_2_io_outputs_2_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_4     (streamDemux_2_io_outputs_2_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_5     (streamDemux_2_io_outputs_2_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_6     (streamDemux_2_io_outputs_2_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_7     (streamDemux_2_io_outputs_2_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_8     (streamDemux_2_io_outputs_2_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_9     (streamDemux_2_io_outputs_2_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_2_payload_0_0_2_10    (streamDemux_2_io_outputs_2_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_11    (streamDemux_2_io_outputs_2_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_12    (streamDemux_2_io_outputs_2_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_13    (streamDemux_2_io_outputs_2_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_14    (streamDemux_2_io_outputs_2_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_2_payload_0_0_2_15    (streamDemux_2_io_outputs_2_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_0     (streamDemux_2_io_outputs_2_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_1     (streamDemux_2_io_outputs_2_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_2     (streamDemux_2_io_outputs_2_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_3     (streamDemux_2_io_outputs_2_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_4     (streamDemux_2_io_outputs_2_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_5     (streamDemux_2_io_outputs_2_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_6     (streamDemux_2_io_outputs_2_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_7     (streamDemux_2_io_outputs_2_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_8     (streamDemux_2_io_outputs_2_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_9     (streamDemux_2_io_outputs_2_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_2_payload_0_1_0_10    (streamDemux_2_io_outputs_2_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_11    (streamDemux_2_io_outputs_2_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_12    (streamDemux_2_io_outputs_2_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_13    (streamDemux_2_io_outputs_2_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_14    (streamDemux_2_io_outputs_2_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_2_payload_0_1_0_15    (streamDemux_2_io_outputs_2_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_0     (streamDemux_2_io_outputs_2_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_1     (streamDemux_2_io_outputs_2_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_2     (streamDemux_2_io_outputs_2_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_3     (streamDemux_2_io_outputs_2_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_4     (streamDemux_2_io_outputs_2_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_5     (streamDemux_2_io_outputs_2_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_6     (streamDemux_2_io_outputs_2_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_7     (streamDemux_2_io_outputs_2_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_8     (streamDemux_2_io_outputs_2_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_9     (streamDemux_2_io_outputs_2_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_2_payload_0_1_1_10    (streamDemux_2_io_outputs_2_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_11    (streamDemux_2_io_outputs_2_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_12    (streamDemux_2_io_outputs_2_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_13    (streamDemux_2_io_outputs_2_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_14    (streamDemux_2_io_outputs_2_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_2_payload_0_1_1_15    (streamDemux_2_io_outputs_2_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_0     (streamDemux_2_io_outputs_2_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_1     (streamDemux_2_io_outputs_2_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_2     (streamDemux_2_io_outputs_2_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_3     (streamDemux_2_io_outputs_2_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_4     (streamDemux_2_io_outputs_2_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_5     (streamDemux_2_io_outputs_2_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_6     (streamDemux_2_io_outputs_2_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_7     (streamDemux_2_io_outputs_2_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_8     (streamDemux_2_io_outputs_2_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_9     (streamDemux_2_io_outputs_2_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_2_payload_0_1_2_10    (streamDemux_2_io_outputs_2_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_11    (streamDemux_2_io_outputs_2_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_12    (streamDemux_2_io_outputs_2_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_13    (streamDemux_2_io_outputs_2_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_14    (streamDemux_2_io_outputs_2_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_2_payload_0_1_2_15    (streamDemux_2_io_outputs_2_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_0     (streamDemux_2_io_outputs_2_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_1     (streamDemux_2_io_outputs_2_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_2     (streamDemux_2_io_outputs_2_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_3     (streamDemux_2_io_outputs_2_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_4     (streamDemux_2_io_outputs_2_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_5     (streamDemux_2_io_outputs_2_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_6     (streamDemux_2_io_outputs_2_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_7     (streamDemux_2_io_outputs_2_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_8     (streamDemux_2_io_outputs_2_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_9     (streamDemux_2_io_outputs_2_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_2_payload_0_2_0_10    (streamDemux_2_io_outputs_2_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_11    (streamDemux_2_io_outputs_2_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_12    (streamDemux_2_io_outputs_2_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_13    (streamDemux_2_io_outputs_2_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_14    (streamDemux_2_io_outputs_2_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_2_payload_0_2_0_15    (streamDemux_2_io_outputs_2_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_0     (streamDemux_2_io_outputs_2_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_1     (streamDemux_2_io_outputs_2_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_2     (streamDemux_2_io_outputs_2_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_3     (streamDemux_2_io_outputs_2_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_4     (streamDemux_2_io_outputs_2_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_5     (streamDemux_2_io_outputs_2_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_6     (streamDemux_2_io_outputs_2_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_7     (streamDemux_2_io_outputs_2_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_8     (streamDemux_2_io_outputs_2_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_9     (streamDemux_2_io_outputs_2_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_2_payload_0_2_1_10    (streamDemux_2_io_outputs_2_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_11    (streamDemux_2_io_outputs_2_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_12    (streamDemux_2_io_outputs_2_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_13    (streamDemux_2_io_outputs_2_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_14    (streamDemux_2_io_outputs_2_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_2_payload_0_2_1_15    (streamDemux_2_io_outputs_2_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_0     (streamDemux_2_io_outputs_2_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_1     (streamDemux_2_io_outputs_2_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_2     (streamDemux_2_io_outputs_2_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_3     (streamDemux_2_io_outputs_2_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_4     (streamDemux_2_io_outputs_2_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_5     (streamDemux_2_io_outputs_2_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_6     (streamDemux_2_io_outputs_2_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_7     (streamDemux_2_io_outputs_2_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_8     (streamDemux_2_io_outputs_2_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_9     (streamDemux_2_io_outputs_2_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_2_payload_0_2_2_10    (streamDemux_2_io_outputs_2_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_11    (streamDemux_2_io_outputs_2_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_12    (streamDemux_2_io_outputs_2_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_13    (streamDemux_2_io_outputs_2_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_14    (streamDemux_2_io_outputs_2_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_2_payload_0_2_2_15    (streamDemux_2_io_outputs_2_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_0     (streamDemux_2_io_outputs_2_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_1     (streamDemux_2_io_outputs_2_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_2     (streamDemux_2_io_outputs_2_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_3     (streamDemux_2_io_outputs_2_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_4     (streamDemux_2_io_outputs_2_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_5     (streamDemux_2_io_outputs_2_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_6     (streamDemux_2_io_outputs_2_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_7     (streamDemux_2_io_outputs_2_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_8     (streamDemux_2_io_outputs_2_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_9     (streamDemux_2_io_outputs_2_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_2_payload_1_0_0_10    (streamDemux_2_io_outputs_2_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_11    (streamDemux_2_io_outputs_2_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_12    (streamDemux_2_io_outputs_2_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_13    (streamDemux_2_io_outputs_2_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_14    (streamDemux_2_io_outputs_2_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_2_payload_1_0_0_15    (streamDemux_2_io_outputs_2_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_0     (streamDemux_2_io_outputs_2_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_1     (streamDemux_2_io_outputs_2_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_2     (streamDemux_2_io_outputs_2_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_3     (streamDemux_2_io_outputs_2_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_4     (streamDemux_2_io_outputs_2_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_5     (streamDemux_2_io_outputs_2_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_6     (streamDemux_2_io_outputs_2_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_7     (streamDemux_2_io_outputs_2_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_8     (streamDemux_2_io_outputs_2_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_9     (streamDemux_2_io_outputs_2_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_2_payload_1_0_1_10    (streamDemux_2_io_outputs_2_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_11    (streamDemux_2_io_outputs_2_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_12    (streamDemux_2_io_outputs_2_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_13    (streamDemux_2_io_outputs_2_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_14    (streamDemux_2_io_outputs_2_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_2_payload_1_0_1_15    (streamDemux_2_io_outputs_2_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_0     (streamDemux_2_io_outputs_2_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_1     (streamDemux_2_io_outputs_2_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_2     (streamDemux_2_io_outputs_2_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_3     (streamDemux_2_io_outputs_2_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_4     (streamDemux_2_io_outputs_2_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_5     (streamDemux_2_io_outputs_2_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_6     (streamDemux_2_io_outputs_2_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_7     (streamDemux_2_io_outputs_2_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_8     (streamDemux_2_io_outputs_2_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_9     (streamDemux_2_io_outputs_2_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_2_payload_1_0_2_10    (streamDemux_2_io_outputs_2_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_11    (streamDemux_2_io_outputs_2_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_12    (streamDemux_2_io_outputs_2_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_13    (streamDemux_2_io_outputs_2_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_14    (streamDemux_2_io_outputs_2_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_2_payload_1_0_2_15    (streamDemux_2_io_outputs_2_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_0     (streamDemux_2_io_outputs_2_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_1     (streamDemux_2_io_outputs_2_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_2     (streamDemux_2_io_outputs_2_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_3     (streamDemux_2_io_outputs_2_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_4     (streamDemux_2_io_outputs_2_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_5     (streamDemux_2_io_outputs_2_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_6     (streamDemux_2_io_outputs_2_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_7     (streamDemux_2_io_outputs_2_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_8     (streamDemux_2_io_outputs_2_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_9     (streamDemux_2_io_outputs_2_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_2_payload_1_1_0_10    (streamDemux_2_io_outputs_2_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_11    (streamDemux_2_io_outputs_2_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_12    (streamDemux_2_io_outputs_2_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_13    (streamDemux_2_io_outputs_2_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_14    (streamDemux_2_io_outputs_2_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_2_payload_1_1_0_15    (streamDemux_2_io_outputs_2_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_0     (streamDemux_2_io_outputs_2_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_1     (streamDemux_2_io_outputs_2_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_2     (streamDemux_2_io_outputs_2_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_3     (streamDemux_2_io_outputs_2_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_4     (streamDemux_2_io_outputs_2_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_5     (streamDemux_2_io_outputs_2_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_6     (streamDemux_2_io_outputs_2_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_7     (streamDemux_2_io_outputs_2_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_8     (streamDemux_2_io_outputs_2_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_9     (streamDemux_2_io_outputs_2_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_2_payload_1_1_1_10    (streamDemux_2_io_outputs_2_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_11    (streamDemux_2_io_outputs_2_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_12    (streamDemux_2_io_outputs_2_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_13    (streamDemux_2_io_outputs_2_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_14    (streamDemux_2_io_outputs_2_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_2_payload_1_1_1_15    (streamDemux_2_io_outputs_2_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_0     (streamDemux_2_io_outputs_2_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_1     (streamDemux_2_io_outputs_2_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_2     (streamDemux_2_io_outputs_2_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_3     (streamDemux_2_io_outputs_2_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_4     (streamDemux_2_io_outputs_2_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_5     (streamDemux_2_io_outputs_2_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_6     (streamDemux_2_io_outputs_2_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_7     (streamDemux_2_io_outputs_2_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_8     (streamDemux_2_io_outputs_2_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_9     (streamDemux_2_io_outputs_2_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_2_payload_1_1_2_10    (streamDemux_2_io_outputs_2_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_11    (streamDemux_2_io_outputs_2_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_12    (streamDemux_2_io_outputs_2_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_13    (streamDemux_2_io_outputs_2_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_14    (streamDemux_2_io_outputs_2_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_2_payload_1_1_2_15    (streamDemux_2_io_outputs_2_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_0     (streamDemux_2_io_outputs_2_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_1     (streamDemux_2_io_outputs_2_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_2     (streamDemux_2_io_outputs_2_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_3     (streamDemux_2_io_outputs_2_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_4     (streamDemux_2_io_outputs_2_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_5     (streamDemux_2_io_outputs_2_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_6     (streamDemux_2_io_outputs_2_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_7     (streamDemux_2_io_outputs_2_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_8     (streamDemux_2_io_outputs_2_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_9     (streamDemux_2_io_outputs_2_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_2_payload_1_2_0_10    (streamDemux_2_io_outputs_2_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_11    (streamDemux_2_io_outputs_2_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_12    (streamDemux_2_io_outputs_2_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_13    (streamDemux_2_io_outputs_2_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_14    (streamDemux_2_io_outputs_2_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_2_payload_1_2_0_15    (streamDemux_2_io_outputs_2_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_0     (streamDemux_2_io_outputs_2_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_1     (streamDemux_2_io_outputs_2_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_2     (streamDemux_2_io_outputs_2_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_3     (streamDemux_2_io_outputs_2_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_4     (streamDemux_2_io_outputs_2_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_5     (streamDemux_2_io_outputs_2_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_6     (streamDemux_2_io_outputs_2_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_7     (streamDemux_2_io_outputs_2_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_8     (streamDemux_2_io_outputs_2_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_9     (streamDemux_2_io_outputs_2_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_2_payload_1_2_1_10    (streamDemux_2_io_outputs_2_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_11    (streamDemux_2_io_outputs_2_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_12    (streamDemux_2_io_outputs_2_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_13    (streamDemux_2_io_outputs_2_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_14    (streamDemux_2_io_outputs_2_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_2_payload_1_2_1_15    (streamDemux_2_io_outputs_2_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_0     (streamDemux_2_io_outputs_2_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_1     (streamDemux_2_io_outputs_2_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_2     (streamDemux_2_io_outputs_2_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_3     (streamDemux_2_io_outputs_2_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_4     (streamDemux_2_io_outputs_2_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_5     (streamDemux_2_io_outputs_2_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_6     (streamDemux_2_io_outputs_2_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_7     (streamDemux_2_io_outputs_2_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_8     (streamDemux_2_io_outputs_2_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_9     (streamDemux_2_io_outputs_2_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_2_payload_1_2_2_10    (streamDemux_2_io_outputs_2_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_11    (streamDemux_2_io_outputs_2_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_12    (streamDemux_2_io_outputs_2_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_13    (streamDemux_2_io_outputs_2_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_14    (streamDemux_2_io_outputs_2_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_2_payload_1_2_2_15    (streamDemux_2_io_outputs_2_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_3_valid               (streamDemux_2_io_outputs_3_valid                  ), //o
    .io_outputs_3_ready               (weightFifo_3_push_ready                           ), //i
    .io_outputs_3_payload_0_0_0_0     (streamDemux_2_io_outputs_3_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_1     (streamDemux_2_io_outputs_3_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_2     (streamDemux_2_io_outputs_3_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_3     (streamDemux_2_io_outputs_3_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_4     (streamDemux_2_io_outputs_3_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_5     (streamDemux_2_io_outputs_3_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_6     (streamDemux_2_io_outputs_3_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_7     (streamDemux_2_io_outputs_3_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_8     (streamDemux_2_io_outputs_3_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_9     (streamDemux_2_io_outputs_3_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_3_payload_0_0_0_10    (streamDemux_2_io_outputs_3_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_3_payload_0_0_0_11    (streamDemux_2_io_outputs_3_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_3_payload_0_0_0_12    (streamDemux_2_io_outputs_3_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_3_payload_0_0_0_13    (streamDemux_2_io_outputs_3_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_3_payload_0_0_0_14    (streamDemux_2_io_outputs_3_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_3_payload_0_0_0_15    (streamDemux_2_io_outputs_3_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_0     (streamDemux_2_io_outputs_3_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_1     (streamDemux_2_io_outputs_3_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_2     (streamDemux_2_io_outputs_3_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_3     (streamDemux_2_io_outputs_3_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_4     (streamDemux_2_io_outputs_3_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_5     (streamDemux_2_io_outputs_3_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_6     (streamDemux_2_io_outputs_3_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_7     (streamDemux_2_io_outputs_3_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_8     (streamDemux_2_io_outputs_3_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_9     (streamDemux_2_io_outputs_3_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_3_payload_0_0_1_10    (streamDemux_2_io_outputs_3_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_11    (streamDemux_2_io_outputs_3_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_12    (streamDemux_2_io_outputs_3_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_13    (streamDemux_2_io_outputs_3_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_14    (streamDemux_2_io_outputs_3_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_3_payload_0_0_1_15    (streamDemux_2_io_outputs_3_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_0     (streamDemux_2_io_outputs_3_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_1     (streamDemux_2_io_outputs_3_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_2     (streamDemux_2_io_outputs_3_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_3     (streamDemux_2_io_outputs_3_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_4     (streamDemux_2_io_outputs_3_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_5     (streamDemux_2_io_outputs_3_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_6     (streamDemux_2_io_outputs_3_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_7     (streamDemux_2_io_outputs_3_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_8     (streamDemux_2_io_outputs_3_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_9     (streamDemux_2_io_outputs_3_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_3_payload_0_0_2_10    (streamDemux_2_io_outputs_3_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_11    (streamDemux_2_io_outputs_3_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_12    (streamDemux_2_io_outputs_3_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_13    (streamDemux_2_io_outputs_3_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_14    (streamDemux_2_io_outputs_3_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_3_payload_0_0_2_15    (streamDemux_2_io_outputs_3_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_0     (streamDemux_2_io_outputs_3_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_1     (streamDemux_2_io_outputs_3_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_2     (streamDemux_2_io_outputs_3_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_3     (streamDemux_2_io_outputs_3_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_4     (streamDemux_2_io_outputs_3_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_5     (streamDemux_2_io_outputs_3_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_6     (streamDemux_2_io_outputs_3_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_7     (streamDemux_2_io_outputs_3_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_8     (streamDemux_2_io_outputs_3_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_9     (streamDemux_2_io_outputs_3_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_3_payload_0_1_0_10    (streamDemux_2_io_outputs_3_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_11    (streamDemux_2_io_outputs_3_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_12    (streamDemux_2_io_outputs_3_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_13    (streamDemux_2_io_outputs_3_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_14    (streamDemux_2_io_outputs_3_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_3_payload_0_1_0_15    (streamDemux_2_io_outputs_3_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_0     (streamDemux_2_io_outputs_3_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_1     (streamDemux_2_io_outputs_3_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_2     (streamDemux_2_io_outputs_3_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_3     (streamDemux_2_io_outputs_3_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_4     (streamDemux_2_io_outputs_3_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_5     (streamDemux_2_io_outputs_3_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_6     (streamDemux_2_io_outputs_3_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_7     (streamDemux_2_io_outputs_3_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_8     (streamDemux_2_io_outputs_3_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_9     (streamDemux_2_io_outputs_3_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_3_payload_0_1_1_10    (streamDemux_2_io_outputs_3_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_11    (streamDemux_2_io_outputs_3_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_12    (streamDemux_2_io_outputs_3_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_13    (streamDemux_2_io_outputs_3_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_14    (streamDemux_2_io_outputs_3_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_3_payload_0_1_1_15    (streamDemux_2_io_outputs_3_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_0     (streamDemux_2_io_outputs_3_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_1     (streamDemux_2_io_outputs_3_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_2     (streamDemux_2_io_outputs_3_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_3     (streamDemux_2_io_outputs_3_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_4     (streamDemux_2_io_outputs_3_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_5     (streamDemux_2_io_outputs_3_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_6     (streamDemux_2_io_outputs_3_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_7     (streamDemux_2_io_outputs_3_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_8     (streamDemux_2_io_outputs_3_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_9     (streamDemux_2_io_outputs_3_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_3_payload_0_1_2_10    (streamDemux_2_io_outputs_3_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_11    (streamDemux_2_io_outputs_3_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_12    (streamDemux_2_io_outputs_3_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_13    (streamDemux_2_io_outputs_3_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_14    (streamDemux_2_io_outputs_3_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_3_payload_0_1_2_15    (streamDemux_2_io_outputs_3_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_0     (streamDemux_2_io_outputs_3_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_1     (streamDemux_2_io_outputs_3_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_2     (streamDemux_2_io_outputs_3_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_3     (streamDemux_2_io_outputs_3_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_4     (streamDemux_2_io_outputs_3_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_5     (streamDemux_2_io_outputs_3_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_6     (streamDemux_2_io_outputs_3_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_7     (streamDemux_2_io_outputs_3_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_8     (streamDemux_2_io_outputs_3_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_9     (streamDemux_2_io_outputs_3_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_3_payload_0_2_0_10    (streamDemux_2_io_outputs_3_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_11    (streamDemux_2_io_outputs_3_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_12    (streamDemux_2_io_outputs_3_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_13    (streamDemux_2_io_outputs_3_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_14    (streamDemux_2_io_outputs_3_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_3_payload_0_2_0_15    (streamDemux_2_io_outputs_3_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_0     (streamDemux_2_io_outputs_3_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_1     (streamDemux_2_io_outputs_3_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_2     (streamDemux_2_io_outputs_3_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_3     (streamDemux_2_io_outputs_3_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_4     (streamDemux_2_io_outputs_3_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_5     (streamDemux_2_io_outputs_3_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_6     (streamDemux_2_io_outputs_3_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_7     (streamDemux_2_io_outputs_3_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_8     (streamDemux_2_io_outputs_3_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_9     (streamDemux_2_io_outputs_3_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_3_payload_0_2_1_10    (streamDemux_2_io_outputs_3_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_11    (streamDemux_2_io_outputs_3_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_12    (streamDemux_2_io_outputs_3_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_13    (streamDemux_2_io_outputs_3_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_14    (streamDemux_2_io_outputs_3_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_3_payload_0_2_1_15    (streamDemux_2_io_outputs_3_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_0     (streamDemux_2_io_outputs_3_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_1     (streamDemux_2_io_outputs_3_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_2     (streamDemux_2_io_outputs_3_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_3     (streamDemux_2_io_outputs_3_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_4     (streamDemux_2_io_outputs_3_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_5     (streamDemux_2_io_outputs_3_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_6     (streamDemux_2_io_outputs_3_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_7     (streamDemux_2_io_outputs_3_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_8     (streamDemux_2_io_outputs_3_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_9     (streamDemux_2_io_outputs_3_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_3_payload_0_2_2_10    (streamDemux_2_io_outputs_3_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_11    (streamDemux_2_io_outputs_3_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_12    (streamDemux_2_io_outputs_3_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_13    (streamDemux_2_io_outputs_3_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_14    (streamDemux_2_io_outputs_3_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_3_payload_0_2_2_15    (streamDemux_2_io_outputs_3_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_0     (streamDemux_2_io_outputs_3_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_1     (streamDemux_2_io_outputs_3_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_2     (streamDemux_2_io_outputs_3_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_3     (streamDemux_2_io_outputs_3_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_4     (streamDemux_2_io_outputs_3_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_5     (streamDemux_2_io_outputs_3_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_6     (streamDemux_2_io_outputs_3_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_7     (streamDemux_2_io_outputs_3_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_8     (streamDemux_2_io_outputs_3_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_9     (streamDemux_2_io_outputs_3_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_3_payload_1_0_0_10    (streamDemux_2_io_outputs_3_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_11    (streamDemux_2_io_outputs_3_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_12    (streamDemux_2_io_outputs_3_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_13    (streamDemux_2_io_outputs_3_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_14    (streamDemux_2_io_outputs_3_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_3_payload_1_0_0_15    (streamDemux_2_io_outputs_3_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_0     (streamDemux_2_io_outputs_3_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_1     (streamDemux_2_io_outputs_3_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_2     (streamDemux_2_io_outputs_3_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_3     (streamDemux_2_io_outputs_3_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_4     (streamDemux_2_io_outputs_3_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_5     (streamDemux_2_io_outputs_3_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_6     (streamDemux_2_io_outputs_3_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_7     (streamDemux_2_io_outputs_3_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_8     (streamDemux_2_io_outputs_3_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_9     (streamDemux_2_io_outputs_3_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_3_payload_1_0_1_10    (streamDemux_2_io_outputs_3_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_11    (streamDemux_2_io_outputs_3_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_12    (streamDemux_2_io_outputs_3_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_13    (streamDemux_2_io_outputs_3_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_14    (streamDemux_2_io_outputs_3_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_3_payload_1_0_1_15    (streamDemux_2_io_outputs_3_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_0     (streamDemux_2_io_outputs_3_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_1     (streamDemux_2_io_outputs_3_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_2     (streamDemux_2_io_outputs_3_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_3     (streamDemux_2_io_outputs_3_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_4     (streamDemux_2_io_outputs_3_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_5     (streamDemux_2_io_outputs_3_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_6     (streamDemux_2_io_outputs_3_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_7     (streamDemux_2_io_outputs_3_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_8     (streamDemux_2_io_outputs_3_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_9     (streamDemux_2_io_outputs_3_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_3_payload_1_0_2_10    (streamDemux_2_io_outputs_3_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_11    (streamDemux_2_io_outputs_3_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_12    (streamDemux_2_io_outputs_3_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_13    (streamDemux_2_io_outputs_3_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_14    (streamDemux_2_io_outputs_3_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_3_payload_1_0_2_15    (streamDemux_2_io_outputs_3_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_0     (streamDemux_2_io_outputs_3_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_1     (streamDemux_2_io_outputs_3_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_2     (streamDemux_2_io_outputs_3_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_3     (streamDemux_2_io_outputs_3_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_4     (streamDemux_2_io_outputs_3_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_5     (streamDemux_2_io_outputs_3_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_6     (streamDemux_2_io_outputs_3_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_7     (streamDemux_2_io_outputs_3_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_8     (streamDemux_2_io_outputs_3_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_9     (streamDemux_2_io_outputs_3_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_3_payload_1_1_0_10    (streamDemux_2_io_outputs_3_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_11    (streamDemux_2_io_outputs_3_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_12    (streamDemux_2_io_outputs_3_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_13    (streamDemux_2_io_outputs_3_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_14    (streamDemux_2_io_outputs_3_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_3_payload_1_1_0_15    (streamDemux_2_io_outputs_3_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_0     (streamDemux_2_io_outputs_3_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_1     (streamDemux_2_io_outputs_3_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_2     (streamDemux_2_io_outputs_3_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_3     (streamDemux_2_io_outputs_3_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_4     (streamDemux_2_io_outputs_3_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_5     (streamDemux_2_io_outputs_3_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_6     (streamDemux_2_io_outputs_3_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_7     (streamDemux_2_io_outputs_3_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_8     (streamDemux_2_io_outputs_3_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_9     (streamDemux_2_io_outputs_3_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_3_payload_1_1_1_10    (streamDemux_2_io_outputs_3_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_11    (streamDemux_2_io_outputs_3_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_12    (streamDemux_2_io_outputs_3_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_13    (streamDemux_2_io_outputs_3_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_14    (streamDemux_2_io_outputs_3_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_3_payload_1_1_1_15    (streamDemux_2_io_outputs_3_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_0     (streamDemux_2_io_outputs_3_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_1     (streamDemux_2_io_outputs_3_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_2     (streamDemux_2_io_outputs_3_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_3     (streamDemux_2_io_outputs_3_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_4     (streamDemux_2_io_outputs_3_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_5     (streamDemux_2_io_outputs_3_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_6     (streamDemux_2_io_outputs_3_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_7     (streamDemux_2_io_outputs_3_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_8     (streamDemux_2_io_outputs_3_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_9     (streamDemux_2_io_outputs_3_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_3_payload_1_1_2_10    (streamDemux_2_io_outputs_3_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_11    (streamDemux_2_io_outputs_3_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_12    (streamDemux_2_io_outputs_3_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_13    (streamDemux_2_io_outputs_3_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_14    (streamDemux_2_io_outputs_3_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_3_payload_1_1_2_15    (streamDemux_2_io_outputs_3_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_0     (streamDemux_2_io_outputs_3_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_1     (streamDemux_2_io_outputs_3_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_2     (streamDemux_2_io_outputs_3_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_3     (streamDemux_2_io_outputs_3_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_4     (streamDemux_2_io_outputs_3_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_5     (streamDemux_2_io_outputs_3_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_6     (streamDemux_2_io_outputs_3_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_7     (streamDemux_2_io_outputs_3_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_8     (streamDemux_2_io_outputs_3_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_9     (streamDemux_2_io_outputs_3_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_3_payload_1_2_0_10    (streamDemux_2_io_outputs_3_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_11    (streamDemux_2_io_outputs_3_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_12    (streamDemux_2_io_outputs_3_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_13    (streamDemux_2_io_outputs_3_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_14    (streamDemux_2_io_outputs_3_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_3_payload_1_2_0_15    (streamDemux_2_io_outputs_3_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_0     (streamDemux_2_io_outputs_3_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_1     (streamDemux_2_io_outputs_3_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_2     (streamDemux_2_io_outputs_3_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_3     (streamDemux_2_io_outputs_3_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_4     (streamDemux_2_io_outputs_3_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_5     (streamDemux_2_io_outputs_3_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_6     (streamDemux_2_io_outputs_3_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_7     (streamDemux_2_io_outputs_3_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_8     (streamDemux_2_io_outputs_3_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_9     (streamDemux_2_io_outputs_3_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_3_payload_1_2_1_10    (streamDemux_2_io_outputs_3_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_11    (streamDemux_2_io_outputs_3_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_12    (streamDemux_2_io_outputs_3_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_13    (streamDemux_2_io_outputs_3_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_14    (streamDemux_2_io_outputs_3_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_3_payload_1_2_1_15    (streamDemux_2_io_outputs_3_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_0     (streamDemux_2_io_outputs_3_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_1     (streamDemux_2_io_outputs_3_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_2     (streamDemux_2_io_outputs_3_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_3     (streamDemux_2_io_outputs_3_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_4     (streamDemux_2_io_outputs_3_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_5     (streamDemux_2_io_outputs_3_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_6     (streamDemux_2_io_outputs_3_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_7     (streamDemux_2_io_outputs_3_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_8     (streamDemux_2_io_outputs_3_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_9     (streamDemux_2_io_outputs_3_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_3_payload_1_2_2_10    (streamDemux_2_io_outputs_3_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_11    (streamDemux_2_io_outputs_3_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_12    (streamDemux_2_io_outputs_3_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_13    (streamDemux_2_io_outputs_3_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_14    (streamDemux_2_io_outputs_3_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_3_payload_1_2_2_15    (streamDemux_2_io_outputs_3_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_4_valid               (streamDemux_2_io_outputs_4_valid                  ), //o
    .io_outputs_4_ready               (weightFifo_4_push_ready                           ), //i
    .io_outputs_4_payload_0_0_0_0     (streamDemux_2_io_outputs_4_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_1     (streamDemux_2_io_outputs_4_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_2     (streamDemux_2_io_outputs_4_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_3     (streamDemux_2_io_outputs_4_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_4     (streamDemux_2_io_outputs_4_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_5     (streamDemux_2_io_outputs_4_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_6     (streamDemux_2_io_outputs_4_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_7     (streamDemux_2_io_outputs_4_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_8     (streamDemux_2_io_outputs_4_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_9     (streamDemux_2_io_outputs_4_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_4_payload_0_0_0_10    (streamDemux_2_io_outputs_4_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_4_payload_0_0_0_11    (streamDemux_2_io_outputs_4_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_4_payload_0_0_0_12    (streamDemux_2_io_outputs_4_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_4_payload_0_0_0_13    (streamDemux_2_io_outputs_4_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_4_payload_0_0_0_14    (streamDemux_2_io_outputs_4_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_4_payload_0_0_0_15    (streamDemux_2_io_outputs_4_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_0     (streamDemux_2_io_outputs_4_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_1     (streamDemux_2_io_outputs_4_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_2     (streamDemux_2_io_outputs_4_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_3     (streamDemux_2_io_outputs_4_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_4     (streamDemux_2_io_outputs_4_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_5     (streamDemux_2_io_outputs_4_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_6     (streamDemux_2_io_outputs_4_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_7     (streamDemux_2_io_outputs_4_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_8     (streamDemux_2_io_outputs_4_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_9     (streamDemux_2_io_outputs_4_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_4_payload_0_0_1_10    (streamDemux_2_io_outputs_4_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_11    (streamDemux_2_io_outputs_4_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_12    (streamDemux_2_io_outputs_4_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_13    (streamDemux_2_io_outputs_4_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_14    (streamDemux_2_io_outputs_4_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_4_payload_0_0_1_15    (streamDemux_2_io_outputs_4_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_0     (streamDemux_2_io_outputs_4_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_1     (streamDemux_2_io_outputs_4_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_2     (streamDemux_2_io_outputs_4_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_3     (streamDemux_2_io_outputs_4_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_4     (streamDemux_2_io_outputs_4_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_5     (streamDemux_2_io_outputs_4_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_6     (streamDemux_2_io_outputs_4_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_7     (streamDemux_2_io_outputs_4_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_8     (streamDemux_2_io_outputs_4_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_9     (streamDemux_2_io_outputs_4_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_4_payload_0_0_2_10    (streamDemux_2_io_outputs_4_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_11    (streamDemux_2_io_outputs_4_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_12    (streamDemux_2_io_outputs_4_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_13    (streamDemux_2_io_outputs_4_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_14    (streamDemux_2_io_outputs_4_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_4_payload_0_0_2_15    (streamDemux_2_io_outputs_4_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_0     (streamDemux_2_io_outputs_4_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_1     (streamDemux_2_io_outputs_4_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_2     (streamDemux_2_io_outputs_4_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_3     (streamDemux_2_io_outputs_4_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_4     (streamDemux_2_io_outputs_4_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_5     (streamDemux_2_io_outputs_4_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_6     (streamDemux_2_io_outputs_4_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_7     (streamDemux_2_io_outputs_4_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_8     (streamDemux_2_io_outputs_4_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_9     (streamDemux_2_io_outputs_4_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_4_payload_0_1_0_10    (streamDemux_2_io_outputs_4_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_11    (streamDemux_2_io_outputs_4_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_12    (streamDemux_2_io_outputs_4_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_13    (streamDemux_2_io_outputs_4_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_14    (streamDemux_2_io_outputs_4_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_4_payload_0_1_0_15    (streamDemux_2_io_outputs_4_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_0     (streamDemux_2_io_outputs_4_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_1     (streamDemux_2_io_outputs_4_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_2     (streamDemux_2_io_outputs_4_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_3     (streamDemux_2_io_outputs_4_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_4     (streamDemux_2_io_outputs_4_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_5     (streamDemux_2_io_outputs_4_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_6     (streamDemux_2_io_outputs_4_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_7     (streamDemux_2_io_outputs_4_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_8     (streamDemux_2_io_outputs_4_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_9     (streamDemux_2_io_outputs_4_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_4_payload_0_1_1_10    (streamDemux_2_io_outputs_4_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_11    (streamDemux_2_io_outputs_4_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_12    (streamDemux_2_io_outputs_4_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_13    (streamDemux_2_io_outputs_4_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_14    (streamDemux_2_io_outputs_4_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_4_payload_0_1_1_15    (streamDemux_2_io_outputs_4_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_0     (streamDemux_2_io_outputs_4_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_1     (streamDemux_2_io_outputs_4_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_2     (streamDemux_2_io_outputs_4_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_3     (streamDemux_2_io_outputs_4_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_4     (streamDemux_2_io_outputs_4_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_5     (streamDemux_2_io_outputs_4_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_6     (streamDemux_2_io_outputs_4_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_7     (streamDemux_2_io_outputs_4_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_8     (streamDemux_2_io_outputs_4_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_9     (streamDemux_2_io_outputs_4_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_4_payload_0_1_2_10    (streamDemux_2_io_outputs_4_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_11    (streamDemux_2_io_outputs_4_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_12    (streamDemux_2_io_outputs_4_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_13    (streamDemux_2_io_outputs_4_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_14    (streamDemux_2_io_outputs_4_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_4_payload_0_1_2_15    (streamDemux_2_io_outputs_4_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_0     (streamDemux_2_io_outputs_4_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_1     (streamDemux_2_io_outputs_4_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_2     (streamDemux_2_io_outputs_4_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_3     (streamDemux_2_io_outputs_4_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_4     (streamDemux_2_io_outputs_4_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_5     (streamDemux_2_io_outputs_4_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_6     (streamDemux_2_io_outputs_4_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_7     (streamDemux_2_io_outputs_4_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_8     (streamDemux_2_io_outputs_4_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_9     (streamDemux_2_io_outputs_4_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_4_payload_0_2_0_10    (streamDemux_2_io_outputs_4_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_11    (streamDemux_2_io_outputs_4_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_12    (streamDemux_2_io_outputs_4_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_13    (streamDemux_2_io_outputs_4_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_14    (streamDemux_2_io_outputs_4_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_4_payload_0_2_0_15    (streamDemux_2_io_outputs_4_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_0     (streamDemux_2_io_outputs_4_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_1     (streamDemux_2_io_outputs_4_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_2     (streamDemux_2_io_outputs_4_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_3     (streamDemux_2_io_outputs_4_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_4     (streamDemux_2_io_outputs_4_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_5     (streamDemux_2_io_outputs_4_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_6     (streamDemux_2_io_outputs_4_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_7     (streamDemux_2_io_outputs_4_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_8     (streamDemux_2_io_outputs_4_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_9     (streamDemux_2_io_outputs_4_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_4_payload_0_2_1_10    (streamDemux_2_io_outputs_4_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_11    (streamDemux_2_io_outputs_4_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_12    (streamDemux_2_io_outputs_4_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_13    (streamDemux_2_io_outputs_4_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_14    (streamDemux_2_io_outputs_4_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_4_payload_0_2_1_15    (streamDemux_2_io_outputs_4_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_0     (streamDemux_2_io_outputs_4_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_1     (streamDemux_2_io_outputs_4_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_2     (streamDemux_2_io_outputs_4_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_3     (streamDemux_2_io_outputs_4_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_4     (streamDemux_2_io_outputs_4_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_5     (streamDemux_2_io_outputs_4_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_6     (streamDemux_2_io_outputs_4_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_7     (streamDemux_2_io_outputs_4_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_8     (streamDemux_2_io_outputs_4_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_9     (streamDemux_2_io_outputs_4_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_4_payload_0_2_2_10    (streamDemux_2_io_outputs_4_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_11    (streamDemux_2_io_outputs_4_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_12    (streamDemux_2_io_outputs_4_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_13    (streamDemux_2_io_outputs_4_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_14    (streamDemux_2_io_outputs_4_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_4_payload_0_2_2_15    (streamDemux_2_io_outputs_4_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_0     (streamDemux_2_io_outputs_4_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_1     (streamDemux_2_io_outputs_4_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_2     (streamDemux_2_io_outputs_4_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_3     (streamDemux_2_io_outputs_4_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_4     (streamDemux_2_io_outputs_4_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_5     (streamDemux_2_io_outputs_4_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_6     (streamDemux_2_io_outputs_4_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_7     (streamDemux_2_io_outputs_4_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_8     (streamDemux_2_io_outputs_4_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_9     (streamDemux_2_io_outputs_4_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_4_payload_1_0_0_10    (streamDemux_2_io_outputs_4_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_11    (streamDemux_2_io_outputs_4_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_12    (streamDemux_2_io_outputs_4_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_13    (streamDemux_2_io_outputs_4_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_14    (streamDemux_2_io_outputs_4_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_4_payload_1_0_0_15    (streamDemux_2_io_outputs_4_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_0     (streamDemux_2_io_outputs_4_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_1     (streamDemux_2_io_outputs_4_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_2     (streamDemux_2_io_outputs_4_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_3     (streamDemux_2_io_outputs_4_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_4     (streamDemux_2_io_outputs_4_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_5     (streamDemux_2_io_outputs_4_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_6     (streamDemux_2_io_outputs_4_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_7     (streamDemux_2_io_outputs_4_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_8     (streamDemux_2_io_outputs_4_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_9     (streamDemux_2_io_outputs_4_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_4_payload_1_0_1_10    (streamDemux_2_io_outputs_4_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_11    (streamDemux_2_io_outputs_4_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_12    (streamDemux_2_io_outputs_4_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_13    (streamDemux_2_io_outputs_4_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_14    (streamDemux_2_io_outputs_4_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_4_payload_1_0_1_15    (streamDemux_2_io_outputs_4_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_0     (streamDemux_2_io_outputs_4_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_1     (streamDemux_2_io_outputs_4_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_2     (streamDemux_2_io_outputs_4_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_3     (streamDemux_2_io_outputs_4_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_4     (streamDemux_2_io_outputs_4_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_5     (streamDemux_2_io_outputs_4_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_6     (streamDemux_2_io_outputs_4_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_7     (streamDemux_2_io_outputs_4_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_8     (streamDemux_2_io_outputs_4_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_9     (streamDemux_2_io_outputs_4_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_4_payload_1_0_2_10    (streamDemux_2_io_outputs_4_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_11    (streamDemux_2_io_outputs_4_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_12    (streamDemux_2_io_outputs_4_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_13    (streamDemux_2_io_outputs_4_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_14    (streamDemux_2_io_outputs_4_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_4_payload_1_0_2_15    (streamDemux_2_io_outputs_4_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_0     (streamDemux_2_io_outputs_4_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_1     (streamDemux_2_io_outputs_4_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_2     (streamDemux_2_io_outputs_4_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_3     (streamDemux_2_io_outputs_4_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_4     (streamDemux_2_io_outputs_4_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_5     (streamDemux_2_io_outputs_4_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_6     (streamDemux_2_io_outputs_4_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_7     (streamDemux_2_io_outputs_4_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_8     (streamDemux_2_io_outputs_4_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_9     (streamDemux_2_io_outputs_4_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_4_payload_1_1_0_10    (streamDemux_2_io_outputs_4_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_11    (streamDemux_2_io_outputs_4_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_12    (streamDemux_2_io_outputs_4_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_13    (streamDemux_2_io_outputs_4_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_14    (streamDemux_2_io_outputs_4_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_4_payload_1_1_0_15    (streamDemux_2_io_outputs_4_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_0     (streamDemux_2_io_outputs_4_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_1     (streamDemux_2_io_outputs_4_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_2     (streamDemux_2_io_outputs_4_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_3     (streamDemux_2_io_outputs_4_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_4     (streamDemux_2_io_outputs_4_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_5     (streamDemux_2_io_outputs_4_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_6     (streamDemux_2_io_outputs_4_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_7     (streamDemux_2_io_outputs_4_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_8     (streamDemux_2_io_outputs_4_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_9     (streamDemux_2_io_outputs_4_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_4_payload_1_1_1_10    (streamDemux_2_io_outputs_4_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_11    (streamDemux_2_io_outputs_4_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_12    (streamDemux_2_io_outputs_4_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_13    (streamDemux_2_io_outputs_4_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_14    (streamDemux_2_io_outputs_4_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_4_payload_1_1_1_15    (streamDemux_2_io_outputs_4_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_0     (streamDemux_2_io_outputs_4_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_1     (streamDemux_2_io_outputs_4_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_2     (streamDemux_2_io_outputs_4_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_3     (streamDemux_2_io_outputs_4_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_4     (streamDemux_2_io_outputs_4_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_5     (streamDemux_2_io_outputs_4_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_6     (streamDemux_2_io_outputs_4_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_7     (streamDemux_2_io_outputs_4_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_8     (streamDemux_2_io_outputs_4_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_9     (streamDemux_2_io_outputs_4_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_4_payload_1_1_2_10    (streamDemux_2_io_outputs_4_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_11    (streamDemux_2_io_outputs_4_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_12    (streamDemux_2_io_outputs_4_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_13    (streamDemux_2_io_outputs_4_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_14    (streamDemux_2_io_outputs_4_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_4_payload_1_1_2_15    (streamDemux_2_io_outputs_4_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_0     (streamDemux_2_io_outputs_4_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_1     (streamDemux_2_io_outputs_4_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_2     (streamDemux_2_io_outputs_4_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_3     (streamDemux_2_io_outputs_4_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_4     (streamDemux_2_io_outputs_4_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_5     (streamDemux_2_io_outputs_4_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_6     (streamDemux_2_io_outputs_4_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_7     (streamDemux_2_io_outputs_4_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_8     (streamDemux_2_io_outputs_4_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_9     (streamDemux_2_io_outputs_4_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_4_payload_1_2_0_10    (streamDemux_2_io_outputs_4_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_11    (streamDemux_2_io_outputs_4_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_12    (streamDemux_2_io_outputs_4_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_13    (streamDemux_2_io_outputs_4_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_14    (streamDemux_2_io_outputs_4_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_4_payload_1_2_0_15    (streamDemux_2_io_outputs_4_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_0     (streamDemux_2_io_outputs_4_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_1     (streamDemux_2_io_outputs_4_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_2     (streamDemux_2_io_outputs_4_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_3     (streamDemux_2_io_outputs_4_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_4     (streamDemux_2_io_outputs_4_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_5     (streamDemux_2_io_outputs_4_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_6     (streamDemux_2_io_outputs_4_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_7     (streamDemux_2_io_outputs_4_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_8     (streamDemux_2_io_outputs_4_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_9     (streamDemux_2_io_outputs_4_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_4_payload_1_2_1_10    (streamDemux_2_io_outputs_4_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_11    (streamDemux_2_io_outputs_4_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_12    (streamDemux_2_io_outputs_4_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_13    (streamDemux_2_io_outputs_4_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_14    (streamDemux_2_io_outputs_4_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_4_payload_1_2_1_15    (streamDemux_2_io_outputs_4_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_0     (streamDemux_2_io_outputs_4_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_1     (streamDemux_2_io_outputs_4_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_2     (streamDemux_2_io_outputs_4_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_3     (streamDemux_2_io_outputs_4_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_4     (streamDemux_2_io_outputs_4_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_5     (streamDemux_2_io_outputs_4_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_6     (streamDemux_2_io_outputs_4_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_7     (streamDemux_2_io_outputs_4_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_8     (streamDemux_2_io_outputs_4_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_9     (streamDemux_2_io_outputs_4_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_4_payload_1_2_2_10    (streamDemux_2_io_outputs_4_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_11    (streamDemux_2_io_outputs_4_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_12    (streamDemux_2_io_outputs_4_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_13    (streamDemux_2_io_outputs_4_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_14    (streamDemux_2_io_outputs_4_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_4_payload_1_2_2_15    (streamDemux_2_io_outputs_4_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_5_valid               (streamDemux_2_io_outputs_5_valid                  ), //o
    .io_outputs_5_ready               (weightFifo_5_push_ready                           ), //i
    .io_outputs_5_payload_0_0_0_0     (streamDemux_2_io_outputs_5_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_1     (streamDemux_2_io_outputs_5_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_2     (streamDemux_2_io_outputs_5_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_3     (streamDemux_2_io_outputs_5_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_4     (streamDemux_2_io_outputs_5_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_5     (streamDemux_2_io_outputs_5_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_6     (streamDemux_2_io_outputs_5_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_7     (streamDemux_2_io_outputs_5_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_8     (streamDemux_2_io_outputs_5_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_9     (streamDemux_2_io_outputs_5_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_5_payload_0_0_0_10    (streamDemux_2_io_outputs_5_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_5_payload_0_0_0_11    (streamDemux_2_io_outputs_5_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_5_payload_0_0_0_12    (streamDemux_2_io_outputs_5_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_5_payload_0_0_0_13    (streamDemux_2_io_outputs_5_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_5_payload_0_0_0_14    (streamDemux_2_io_outputs_5_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_5_payload_0_0_0_15    (streamDemux_2_io_outputs_5_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_0     (streamDemux_2_io_outputs_5_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_1     (streamDemux_2_io_outputs_5_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_2     (streamDemux_2_io_outputs_5_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_3     (streamDemux_2_io_outputs_5_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_4     (streamDemux_2_io_outputs_5_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_5     (streamDemux_2_io_outputs_5_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_6     (streamDemux_2_io_outputs_5_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_7     (streamDemux_2_io_outputs_5_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_8     (streamDemux_2_io_outputs_5_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_9     (streamDemux_2_io_outputs_5_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_5_payload_0_0_1_10    (streamDemux_2_io_outputs_5_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_11    (streamDemux_2_io_outputs_5_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_12    (streamDemux_2_io_outputs_5_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_13    (streamDemux_2_io_outputs_5_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_14    (streamDemux_2_io_outputs_5_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_5_payload_0_0_1_15    (streamDemux_2_io_outputs_5_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_0     (streamDemux_2_io_outputs_5_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_1     (streamDemux_2_io_outputs_5_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_2     (streamDemux_2_io_outputs_5_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_3     (streamDemux_2_io_outputs_5_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_4     (streamDemux_2_io_outputs_5_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_5     (streamDemux_2_io_outputs_5_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_6     (streamDemux_2_io_outputs_5_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_7     (streamDemux_2_io_outputs_5_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_8     (streamDemux_2_io_outputs_5_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_9     (streamDemux_2_io_outputs_5_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_5_payload_0_0_2_10    (streamDemux_2_io_outputs_5_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_11    (streamDemux_2_io_outputs_5_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_12    (streamDemux_2_io_outputs_5_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_13    (streamDemux_2_io_outputs_5_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_14    (streamDemux_2_io_outputs_5_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_5_payload_0_0_2_15    (streamDemux_2_io_outputs_5_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_0     (streamDemux_2_io_outputs_5_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_1     (streamDemux_2_io_outputs_5_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_2     (streamDemux_2_io_outputs_5_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_3     (streamDemux_2_io_outputs_5_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_4     (streamDemux_2_io_outputs_5_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_5     (streamDemux_2_io_outputs_5_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_6     (streamDemux_2_io_outputs_5_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_7     (streamDemux_2_io_outputs_5_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_8     (streamDemux_2_io_outputs_5_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_9     (streamDemux_2_io_outputs_5_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_5_payload_0_1_0_10    (streamDemux_2_io_outputs_5_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_11    (streamDemux_2_io_outputs_5_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_12    (streamDemux_2_io_outputs_5_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_13    (streamDemux_2_io_outputs_5_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_14    (streamDemux_2_io_outputs_5_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_5_payload_0_1_0_15    (streamDemux_2_io_outputs_5_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_0     (streamDemux_2_io_outputs_5_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_1     (streamDemux_2_io_outputs_5_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_2     (streamDemux_2_io_outputs_5_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_3     (streamDemux_2_io_outputs_5_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_4     (streamDemux_2_io_outputs_5_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_5     (streamDemux_2_io_outputs_5_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_6     (streamDemux_2_io_outputs_5_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_7     (streamDemux_2_io_outputs_5_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_8     (streamDemux_2_io_outputs_5_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_9     (streamDemux_2_io_outputs_5_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_5_payload_0_1_1_10    (streamDemux_2_io_outputs_5_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_11    (streamDemux_2_io_outputs_5_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_12    (streamDemux_2_io_outputs_5_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_13    (streamDemux_2_io_outputs_5_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_14    (streamDemux_2_io_outputs_5_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_5_payload_0_1_1_15    (streamDemux_2_io_outputs_5_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_0     (streamDemux_2_io_outputs_5_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_1     (streamDemux_2_io_outputs_5_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_2     (streamDemux_2_io_outputs_5_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_3     (streamDemux_2_io_outputs_5_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_4     (streamDemux_2_io_outputs_5_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_5     (streamDemux_2_io_outputs_5_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_6     (streamDemux_2_io_outputs_5_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_7     (streamDemux_2_io_outputs_5_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_8     (streamDemux_2_io_outputs_5_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_9     (streamDemux_2_io_outputs_5_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_5_payload_0_1_2_10    (streamDemux_2_io_outputs_5_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_11    (streamDemux_2_io_outputs_5_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_12    (streamDemux_2_io_outputs_5_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_13    (streamDemux_2_io_outputs_5_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_14    (streamDemux_2_io_outputs_5_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_5_payload_0_1_2_15    (streamDemux_2_io_outputs_5_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_0     (streamDemux_2_io_outputs_5_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_1     (streamDemux_2_io_outputs_5_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_2     (streamDemux_2_io_outputs_5_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_3     (streamDemux_2_io_outputs_5_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_4     (streamDemux_2_io_outputs_5_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_5     (streamDemux_2_io_outputs_5_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_6     (streamDemux_2_io_outputs_5_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_7     (streamDemux_2_io_outputs_5_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_8     (streamDemux_2_io_outputs_5_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_9     (streamDemux_2_io_outputs_5_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_5_payload_0_2_0_10    (streamDemux_2_io_outputs_5_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_11    (streamDemux_2_io_outputs_5_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_12    (streamDemux_2_io_outputs_5_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_13    (streamDemux_2_io_outputs_5_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_14    (streamDemux_2_io_outputs_5_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_5_payload_0_2_0_15    (streamDemux_2_io_outputs_5_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_0     (streamDemux_2_io_outputs_5_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_1     (streamDemux_2_io_outputs_5_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_2     (streamDemux_2_io_outputs_5_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_3     (streamDemux_2_io_outputs_5_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_4     (streamDemux_2_io_outputs_5_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_5     (streamDemux_2_io_outputs_5_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_6     (streamDemux_2_io_outputs_5_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_7     (streamDemux_2_io_outputs_5_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_8     (streamDemux_2_io_outputs_5_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_9     (streamDemux_2_io_outputs_5_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_5_payload_0_2_1_10    (streamDemux_2_io_outputs_5_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_11    (streamDemux_2_io_outputs_5_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_12    (streamDemux_2_io_outputs_5_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_13    (streamDemux_2_io_outputs_5_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_14    (streamDemux_2_io_outputs_5_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_5_payload_0_2_1_15    (streamDemux_2_io_outputs_5_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_0     (streamDemux_2_io_outputs_5_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_1     (streamDemux_2_io_outputs_5_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_2     (streamDemux_2_io_outputs_5_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_3     (streamDemux_2_io_outputs_5_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_4     (streamDemux_2_io_outputs_5_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_5     (streamDemux_2_io_outputs_5_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_6     (streamDemux_2_io_outputs_5_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_7     (streamDemux_2_io_outputs_5_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_8     (streamDemux_2_io_outputs_5_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_9     (streamDemux_2_io_outputs_5_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_5_payload_0_2_2_10    (streamDemux_2_io_outputs_5_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_11    (streamDemux_2_io_outputs_5_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_12    (streamDemux_2_io_outputs_5_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_13    (streamDemux_2_io_outputs_5_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_14    (streamDemux_2_io_outputs_5_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_5_payload_0_2_2_15    (streamDemux_2_io_outputs_5_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_0     (streamDemux_2_io_outputs_5_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_1     (streamDemux_2_io_outputs_5_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_2     (streamDemux_2_io_outputs_5_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_3     (streamDemux_2_io_outputs_5_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_4     (streamDemux_2_io_outputs_5_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_5     (streamDemux_2_io_outputs_5_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_6     (streamDemux_2_io_outputs_5_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_7     (streamDemux_2_io_outputs_5_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_8     (streamDemux_2_io_outputs_5_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_9     (streamDemux_2_io_outputs_5_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_5_payload_1_0_0_10    (streamDemux_2_io_outputs_5_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_11    (streamDemux_2_io_outputs_5_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_12    (streamDemux_2_io_outputs_5_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_13    (streamDemux_2_io_outputs_5_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_14    (streamDemux_2_io_outputs_5_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_5_payload_1_0_0_15    (streamDemux_2_io_outputs_5_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_0     (streamDemux_2_io_outputs_5_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_1     (streamDemux_2_io_outputs_5_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_2     (streamDemux_2_io_outputs_5_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_3     (streamDemux_2_io_outputs_5_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_4     (streamDemux_2_io_outputs_5_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_5     (streamDemux_2_io_outputs_5_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_6     (streamDemux_2_io_outputs_5_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_7     (streamDemux_2_io_outputs_5_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_8     (streamDemux_2_io_outputs_5_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_9     (streamDemux_2_io_outputs_5_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_5_payload_1_0_1_10    (streamDemux_2_io_outputs_5_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_11    (streamDemux_2_io_outputs_5_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_12    (streamDemux_2_io_outputs_5_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_13    (streamDemux_2_io_outputs_5_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_14    (streamDemux_2_io_outputs_5_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_5_payload_1_0_1_15    (streamDemux_2_io_outputs_5_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_0     (streamDemux_2_io_outputs_5_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_1     (streamDemux_2_io_outputs_5_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_2     (streamDemux_2_io_outputs_5_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_3     (streamDemux_2_io_outputs_5_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_4     (streamDemux_2_io_outputs_5_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_5     (streamDemux_2_io_outputs_5_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_6     (streamDemux_2_io_outputs_5_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_7     (streamDemux_2_io_outputs_5_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_8     (streamDemux_2_io_outputs_5_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_9     (streamDemux_2_io_outputs_5_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_5_payload_1_0_2_10    (streamDemux_2_io_outputs_5_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_11    (streamDemux_2_io_outputs_5_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_12    (streamDemux_2_io_outputs_5_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_13    (streamDemux_2_io_outputs_5_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_14    (streamDemux_2_io_outputs_5_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_5_payload_1_0_2_15    (streamDemux_2_io_outputs_5_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_0     (streamDemux_2_io_outputs_5_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_1     (streamDemux_2_io_outputs_5_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_2     (streamDemux_2_io_outputs_5_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_3     (streamDemux_2_io_outputs_5_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_4     (streamDemux_2_io_outputs_5_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_5     (streamDemux_2_io_outputs_5_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_6     (streamDemux_2_io_outputs_5_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_7     (streamDemux_2_io_outputs_5_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_8     (streamDemux_2_io_outputs_5_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_9     (streamDemux_2_io_outputs_5_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_5_payload_1_1_0_10    (streamDemux_2_io_outputs_5_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_11    (streamDemux_2_io_outputs_5_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_12    (streamDemux_2_io_outputs_5_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_13    (streamDemux_2_io_outputs_5_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_14    (streamDemux_2_io_outputs_5_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_5_payload_1_1_0_15    (streamDemux_2_io_outputs_5_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_0     (streamDemux_2_io_outputs_5_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_1     (streamDemux_2_io_outputs_5_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_2     (streamDemux_2_io_outputs_5_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_3     (streamDemux_2_io_outputs_5_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_4     (streamDemux_2_io_outputs_5_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_5     (streamDemux_2_io_outputs_5_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_6     (streamDemux_2_io_outputs_5_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_7     (streamDemux_2_io_outputs_5_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_8     (streamDemux_2_io_outputs_5_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_9     (streamDemux_2_io_outputs_5_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_5_payload_1_1_1_10    (streamDemux_2_io_outputs_5_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_11    (streamDemux_2_io_outputs_5_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_12    (streamDemux_2_io_outputs_5_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_13    (streamDemux_2_io_outputs_5_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_14    (streamDemux_2_io_outputs_5_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_5_payload_1_1_1_15    (streamDemux_2_io_outputs_5_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_0     (streamDemux_2_io_outputs_5_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_1     (streamDemux_2_io_outputs_5_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_2     (streamDemux_2_io_outputs_5_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_3     (streamDemux_2_io_outputs_5_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_4     (streamDemux_2_io_outputs_5_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_5     (streamDemux_2_io_outputs_5_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_6     (streamDemux_2_io_outputs_5_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_7     (streamDemux_2_io_outputs_5_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_8     (streamDemux_2_io_outputs_5_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_9     (streamDemux_2_io_outputs_5_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_5_payload_1_1_2_10    (streamDemux_2_io_outputs_5_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_11    (streamDemux_2_io_outputs_5_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_12    (streamDemux_2_io_outputs_5_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_13    (streamDemux_2_io_outputs_5_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_14    (streamDemux_2_io_outputs_5_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_5_payload_1_1_2_15    (streamDemux_2_io_outputs_5_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_0     (streamDemux_2_io_outputs_5_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_1     (streamDemux_2_io_outputs_5_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_2     (streamDemux_2_io_outputs_5_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_3     (streamDemux_2_io_outputs_5_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_4     (streamDemux_2_io_outputs_5_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_5     (streamDemux_2_io_outputs_5_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_6     (streamDemux_2_io_outputs_5_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_7     (streamDemux_2_io_outputs_5_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_8     (streamDemux_2_io_outputs_5_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_9     (streamDemux_2_io_outputs_5_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_5_payload_1_2_0_10    (streamDemux_2_io_outputs_5_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_11    (streamDemux_2_io_outputs_5_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_12    (streamDemux_2_io_outputs_5_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_13    (streamDemux_2_io_outputs_5_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_14    (streamDemux_2_io_outputs_5_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_5_payload_1_2_0_15    (streamDemux_2_io_outputs_5_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_0     (streamDemux_2_io_outputs_5_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_1     (streamDemux_2_io_outputs_5_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_2     (streamDemux_2_io_outputs_5_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_3     (streamDemux_2_io_outputs_5_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_4     (streamDemux_2_io_outputs_5_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_5     (streamDemux_2_io_outputs_5_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_6     (streamDemux_2_io_outputs_5_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_7     (streamDemux_2_io_outputs_5_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_8     (streamDemux_2_io_outputs_5_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_9     (streamDemux_2_io_outputs_5_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_5_payload_1_2_1_10    (streamDemux_2_io_outputs_5_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_11    (streamDemux_2_io_outputs_5_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_12    (streamDemux_2_io_outputs_5_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_13    (streamDemux_2_io_outputs_5_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_14    (streamDemux_2_io_outputs_5_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_5_payload_1_2_1_15    (streamDemux_2_io_outputs_5_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_0     (streamDemux_2_io_outputs_5_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_1     (streamDemux_2_io_outputs_5_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_2     (streamDemux_2_io_outputs_5_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_3     (streamDemux_2_io_outputs_5_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_4     (streamDemux_2_io_outputs_5_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_5     (streamDemux_2_io_outputs_5_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_6     (streamDemux_2_io_outputs_5_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_7     (streamDemux_2_io_outputs_5_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_8     (streamDemux_2_io_outputs_5_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_9     (streamDemux_2_io_outputs_5_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_5_payload_1_2_2_10    (streamDemux_2_io_outputs_5_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_11    (streamDemux_2_io_outputs_5_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_12    (streamDemux_2_io_outputs_5_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_13    (streamDemux_2_io_outputs_5_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_14    (streamDemux_2_io_outputs_5_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_5_payload_1_2_2_15    (streamDemux_2_io_outputs_5_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_6_valid               (streamDemux_2_io_outputs_6_valid                  ), //o
    .io_outputs_6_ready               (weightFifo_6_push_ready                           ), //i
    .io_outputs_6_payload_0_0_0_0     (streamDemux_2_io_outputs_6_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_1     (streamDemux_2_io_outputs_6_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_2     (streamDemux_2_io_outputs_6_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_3     (streamDemux_2_io_outputs_6_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_4     (streamDemux_2_io_outputs_6_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_5     (streamDemux_2_io_outputs_6_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_6     (streamDemux_2_io_outputs_6_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_7     (streamDemux_2_io_outputs_6_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_8     (streamDemux_2_io_outputs_6_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_9     (streamDemux_2_io_outputs_6_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_6_payload_0_0_0_10    (streamDemux_2_io_outputs_6_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_6_payload_0_0_0_11    (streamDemux_2_io_outputs_6_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_6_payload_0_0_0_12    (streamDemux_2_io_outputs_6_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_6_payload_0_0_0_13    (streamDemux_2_io_outputs_6_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_6_payload_0_0_0_14    (streamDemux_2_io_outputs_6_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_6_payload_0_0_0_15    (streamDemux_2_io_outputs_6_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_0     (streamDemux_2_io_outputs_6_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_1     (streamDemux_2_io_outputs_6_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_2     (streamDemux_2_io_outputs_6_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_3     (streamDemux_2_io_outputs_6_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_4     (streamDemux_2_io_outputs_6_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_5     (streamDemux_2_io_outputs_6_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_6     (streamDemux_2_io_outputs_6_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_7     (streamDemux_2_io_outputs_6_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_8     (streamDemux_2_io_outputs_6_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_9     (streamDemux_2_io_outputs_6_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_6_payload_0_0_1_10    (streamDemux_2_io_outputs_6_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_11    (streamDemux_2_io_outputs_6_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_12    (streamDemux_2_io_outputs_6_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_13    (streamDemux_2_io_outputs_6_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_14    (streamDemux_2_io_outputs_6_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_6_payload_0_0_1_15    (streamDemux_2_io_outputs_6_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_0     (streamDemux_2_io_outputs_6_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_1     (streamDemux_2_io_outputs_6_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_2     (streamDemux_2_io_outputs_6_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_3     (streamDemux_2_io_outputs_6_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_4     (streamDemux_2_io_outputs_6_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_5     (streamDemux_2_io_outputs_6_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_6     (streamDemux_2_io_outputs_6_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_7     (streamDemux_2_io_outputs_6_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_8     (streamDemux_2_io_outputs_6_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_9     (streamDemux_2_io_outputs_6_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_6_payload_0_0_2_10    (streamDemux_2_io_outputs_6_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_11    (streamDemux_2_io_outputs_6_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_12    (streamDemux_2_io_outputs_6_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_13    (streamDemux_2_io_outputs_6_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_14    (streamDemux_2_io_outputs_6_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_6_payload_0_0_2_15    (streamDemux_2_io_outputs_6_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_0     (streamDemux_2_io_outputs_6_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_1     (streamDemux_2_io_outputs_6_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_2     (streamDemux_2_io_outputs_6_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_3     (streamDemux_2_io_outputs_6_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_4     (streamDemux_2_io_outputs_6_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_5     (streamDemux_2_io_outputs_6_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_6     (streamDemux_2_io_outputs_6_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_7     (streamDemux_2_io_outputs_6_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_8     (streamDemux_2_io_outputs_6_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_9     (streamDemux_2_io_outputs_6_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_6_payload_0_1_0_10    (streamDemux_2_io_outputs_6_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_11    (streamDemux_2_io_outputs_6_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_12    (streamDemux_2_io_outputs_6_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_13    (streamDemux_2_io_outputs_6_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_14    (streamDemux_2_io_outputs_6_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_6_payload_0_1_0_15    (streamDemux_2_io_outputs_6_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_0     (streamDemux_2_io_outputs_6_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_1     (streamDemux_2_io_outputs_6_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_2     (streamDemux_2_io_outputs_6_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_3     (streamDemux_2_io_outputs_6_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_4     (streamDemux_2_io_outputs_6_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_5     (streamDemux_2_io_outputs_6_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_6     (streamDemux_2_io_outputs_6_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_7     (streamDemux_2_io_outputs_6_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_8     (streamDemux_2_io_outputs_6_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_9     (streamDemux_2_io_outputs_6_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_6_payload_0_1_1_10    (streamDemux_2_io_outputs_6_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_11    (streamDemux_2_io_outputs_6_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_12    (streamDemux_2_io_outputs_6_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_13    (streamDemux_2_io_outputs_6_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_14    (streamDemux_2_io_outputs_6_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_6_payload_0_1_1_15    (streamDemux_2_io_outputs_6_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_0     (streamDemux_2_io_outputs_6_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_1     (streamDemux_2_io_outputs_6_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_2     (streamDemux_2_io_outputs_6_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_3     (streamDemux_2_io_outputs_6_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_4     (streamDemux_2_io_outputs_6_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_5     (streamDemux_2_io_outputs_6_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_6     (streamDemux_2_io_outputs_6_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_7     (streamDemux_2_io_outputs_6_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_8     (streamDemux_2_io_outputs_6_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_9     (streamDemux_2_io_outputs_6_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_6_payload_0_1_2_10    (streamDemux_2_io_outputs_6_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_11    (streamDemux_2_io_outputs_6_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_12    (streamDemux_2_io_outputs_6_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_13    (streamDemux_2_io_outputs_6_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_14    (streamDemux_2_io_outputs_6_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_6_payload_0_1_2_15    (streamDemux_2_io_outputs_6_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_0     (streamDemux_2_io_outputs_6_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_1     (streamDemux_2_io_outputs_6_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_2     (streamDemux_2_io_outputs_6_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_3     (streamDemux_2_io_outputs_6_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_4     (streamDemux_2_io_outputs_6_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_5     (streamDemux_2_io_outputs_6_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_6     (streamDemux_2_io_outputs_6_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_7     (streamDemux_2_io_outputs_6_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_8     (streamDemux_2_io_outputs_6_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_9     (streamDemux_2_io_outputs_6_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_6_payload_0_2_0_10    (streamDemux_2_io_outputs_6_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_11    (streamDemux_2_io_outputs_6_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_12    (streamDemux_2_io_outputs_6_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_13    (streamDemux_2_io_outputs_6_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_14    (streamDemux_2_io_outputs_6_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_6_payload_0_2_0_15    (streamDemux_2_io_outputs_6_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_0     (streamDemux_2_io_outputs_6_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_1     (streamDemux_2_io_outputs_6_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_2     (streamDemux_2_io_outputs_6_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_3     (streamDemux_2_io_outputs_6_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_4     (streamDemux_2_io_outputs_6_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_5     (streamDemux_2_io_outputs_6_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_6     (streamDemux_2_io_outputs_6_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_7     (streamDemux_2_io_outputs_6_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_8     (streamDemux_2_io_outputs_6_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_9     (streamDemux_2_io_outputs_6_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_6_payload_0_2_1_10    (streamDemux_2_io_outputs_6_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_11    (streamDemux_2_io_outputs_6_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_12    (streamDemux_2_io_outputs_6_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_13    (streamDemux_2_io_outputs_6_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_14    (streamDemux_2_io_outputs_6_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_6_payload_0_2_1_15    (streamDemux_2_io_outputs_6_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_0     (streamDemux_2_io_outputs_6_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_1     (streamDemux_2_io_outputs_6_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_2     (streamDemux_2_io_outputs_6_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_3     (streamDemux_2_io_outputs_6_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_4     (streamDemux_2_io_outputs_6_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_5     (streamDemux_2_io_outputs_6_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_6     (streamDemux_2_io_outputs_6_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_7     (streamDemux_2_io_outputs_6_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_8     (streamDemux_2_io_outputs_6_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_9     (streamDemux_2_io_outputs_6_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_6_payload_0_2_2_10    (streamDemux_2_io_outputs_6_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_11    (streamDemux_2_io_outputs_6_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_12    (streamDemux_2_io_outputs_6_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_13    (streamDemux_2_io_outputs_6_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_14    (streamDemux_2_io_outputs_6_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_6_payload_0_2_2_15    (streamDemux_2_io_outputs_6_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_0     (streamDemux_2_io_outputs_6_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_1     (streamDemux_2_io_outputs_6_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_2     (streamDemux_2_io_outputs_6_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_3     (streamDemux_2_io_outputs_6_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_4     (streamDemux_2_io_outputs_6_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_5     (streamDemux_2_io_outputs_6_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_6     (streamDemux_2_io_outputs_6_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_7     (streamDemux_2_io_outputs_6_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_8     (streamDemux_2_io_outputs_6_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_9     (streamDemux_2_io_outputs_6_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_6_payload_1_0_0_10    (streamDemux_2_io_outputs_6_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_11    (streamDemux_2_io_outputs_6_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_12    (streamDemux_2_io_outputs_6_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_13    (streamDemux_2_io_outputs_6_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_14    (streamDemux_2_io_outputs_6_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_6_payload_1_0_0_15    (streamDemux_2_io_outputs_6_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_0     (streamDemux_2_io_outputs_6_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_1     (streamDemux_2_io_outputs_6_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_2     (streamDemux_2_io_outputs_6_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_3     (streamDemux_2_io_outputs_6_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_4     (streamDemux_2_io_outputs_6_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_5     (streamDemux_2_io_outputs_6_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_6     (streamDemux_2_io_outputs_6_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_7     (streamDemux_2_io_outputs_6_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_8     (streamDemux_2_io_outputs_6_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_9     (streamDemux_2_io_outputs_6_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_6_payload_1_0_1_10    (streamDemux_2_io_outputs_6_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_11    (streamDemux_2_io_outputs_6_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_12    (streamDemux_2_io_outputs_6_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_13    (streamDemux_2_io_outputs_6_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_14    (streamDemux_2_io_outputs_6_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_6_payload_1_0_1_15    (streamDemux_2_io_outputs_6_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_0     (streamDemux_2_io_outputs_6_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_1     (streamDemux_2_io_outputs_6_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_2     (streamDemux_2_io_outputs_6_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_3     (streamDemux_2_io_outputs_6_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_4     (streamDemux_2_io_outputs_6_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_5     (streamDemux_2_io_outputs_6_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_6     (streamDemux_2_io_outputs_6_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_7     (streamDemux_2_io_outputs_6_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_8     (streamDemux_2_io_outputs_6_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_9     (streamDemux_2_io_outputs_6_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_6_payload_1_0_2_10    (streamDemux_2_io_outputs_6_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_11    (streamDemux_2_io_outputs_6_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_12    (streamDemux_2_io_outputs_6_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_13    (streamDemux_2_io_outputs_6_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_14    (streamDemux_2_io_outputs_6_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_6_payload_1_0_2_15    (streamDemux_2_io_outputs_6_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_0     (streamDemux_2_io_outputs_6_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_1     (streamDemux_2_io_outputs_6_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_2     (streamDemux_2_io_outputs_6_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_3     (streamDemux_2_io_outputs_6_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_4     (streamDemux_2_io_outputs_6_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_5     (streamDemux_2_io_outputs_6_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_6     (streamDemux_2_io_outputs_6_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_7     (streamDemux_2_io_outputs_6_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_8     (streamDemux_2_io_outputs_6_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_9     (streamDemux_2_io_outputs_6_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_6_payload_1_1_0_10    (streamDemux_2_io_outputs_6_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_11    (streamDemux_2_io_outputs_6_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_12    (streamDemux_2_io_outputs_6_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_13    (streamDemux_2_io_outputs_6_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_14    (streamDemux_2_io_outputs_6_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_6_payload_1_1_0_15    (streamDemux_2_io_outputs_6_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_0     (streamDemux_2_io_outputs_6_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_1     (streamDemux_2_io_outputs_6_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_2     (streamDemux_2_io_outputs_6_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_3     (streamDemux_2_io_outputs_6_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_4     (streamDemux_2_io_outputs_6_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_5     (streamDemux_2_io_outputs_6_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_6     (streamDemux_2_io_outputs_6_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_7     (streamDemux_2_io_outputs_6_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_8     (streamDemux_2_io_outputs_6_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_9     (streamDemux_2_io_outputs_6_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_6_payload_1_1_1_10    (streamDemux_2_io_outputs_6_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_11    (streamDemux_2_io_outputs_6_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_12    (streamDemux_2_io_outputs_6_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_13    (streamDemux_2_io_outputs_6_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_14    (streamDemux_2_io_outputs_6_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_6_payload_1_1_1_15    (streamDemux_2_io_outputs_6_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_0     (streamDemux_2_io_outputs_6_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_1     (streamDemux_2_io_outputs_6_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_2     (streamDemux_2_io_outputs_6_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_3     (streamDemux_2_io_outputs_6_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_4     (streamDemux_2_io_outputs_6_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_5     (streamDemux_2_io_outputs_6_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_6     (streamDemux_2_io_outputs_6_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_7     (streamDemux_2_io_outputs_6_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_8     (streamDemux_2_io_outputs_6_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_9     (streamDemux_2_io_outputs_6_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_6_payload_1_1_2_10    (streamDemux_2_io_outputs_6_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_11    (streamDemux_2_io_outputs_6_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_12    (streamDemux_2_io_outputs_6_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_13    (streamDemux_2_io_outputs_6_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_14    (streamDemux_2_io_outputs_6_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_6_payload_1_1_2_15    (streamDemux_2_io_outputs_6_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_0     (streamDemux_2_io_outputs_6_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_1     (streamDemux_2_io_outputs_6_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_2     (streamDemux_2_io_outputs_6_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_3     (streamDemux_2_io_outputs_6_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_4     (streamDemux_2_io_outputs_6_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_5     (streamDemux_2_io_outputs_6_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_6     (streamDemux_2_io_outputs_6_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_7     (streamDemux_2_io_outputs_6_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_8     (streamDemux_2_io_outputs_6_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_9     (streamDemux_2_io_outputs_6_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_6_payload_1_2_0_10    (streamDemux_2_io_outputs_6_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_11    (streamDemux_2_io_outputs_6_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_12    (streamDemux_2_io_outputs_6_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_13    (streamDemux_2_io_outputs_6_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_14    (streamDemux_2_io_outputs_6_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_6_payload_1_2_0_15    (streamDemux_2_io_outputs_6_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_0     (streamDemux_2_io_outputs_6_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_1     (streamDemux_2_io_outputs_6_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_2     (streamDemux_2_io_outputs_6_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_3     (streamDemux_2_io_outputs_6_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_4     (streamDemux_2_io_outputs_6_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_5     (streamDemux_2_io_outputs_6_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_6     (streamDemux_2_io_outputs_6_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_7     (streamDemux_2_io_outputs_6_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_8     (streamDemux_2_io_outputs_6_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_9     (streamDemux_2_io_outputs_6_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_6_payload_1_2_1_10    (streamDemux_2_io_outputs_6_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_11    (streamDemux_2_io_outputs_6_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_12    (streamDemux_2_io_outputs_6_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_13    (streamDemux_2_io_outputs_6_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_14    (streamDemux_2_io_outputs_6_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_6_payload_1_2_1_15    (streamDemux_2_io_outputs_6_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_0     (streamDemux_2_io_outputs_6_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_1     (streamDemux_2_io_outputs_6_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_2     (streamDemux_2_io_outputs_6_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_3     (streamDemux_2_io_outputs_6_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_4     (streamDemux_2_io_outputs_6_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_5     (streamDemux_2_io_outputs_6_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_6     (streamDemux_2_io_outputs_6_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_7     (streamDemux_2_io_outputs_6_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_8     (streamDemux_2_io_outputs_6_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_9     (streamDemux_2_io_outputs_6_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_6_payload_1_2_2_10    (streamDemux_2_io_outputs_6_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_11    (streamDemux_2_io_outputs_6_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_12    (streamDemux_2_io_outputs_6_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_13    (streamDemux_2_io_outputs_6_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_14    (streamDemux_2_io_outputs_6_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_6_payload_1_2_2_15    (streamDemux_2_io_outputs_6_payload_1_2_2_15[7:0]  ), //o
    .io_outputs_7_valid               (streamDemux_2_io_outputs_7_valid                  ), //o
    .io_outputs_7_ready               (weightFifo_7_push_ready                           ), //i
    .io_outputs_7_payload_0_0_0_0     (streamDemux_2_io_outputs_7_payload_0_0_0_0[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_1     (streamDemux_2_io_outputs_7_payload_0_0_0_1[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_2     (streamDemux_2_io_outputs_7_payload_0_0_0_2[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_3     (streamDemux_2_io_outputs_7_payload_0_0_0_3[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_4     (streamDemux_2_io_outputs_7_payload_0_0_0_4[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_5     (streamDemux_2_io_outputs_7_payload_0_0_0_5[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_6     (streamDemux_2_io_outputs_7_payload_0_0_0_6[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_7     (streamDemux_2_io_outputs_7_payload_0_0_0_7[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_8     (streamDemux_2_io_outputs_7_payload_0_0_0_8[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_9     (streamDemux_2_io_outputs_7_payload_0_0_0_9[7:0]   ), //o
    .io_outputs_7_payload_0_0_0_10    (streamDemux_2_io_outputs_7_payload_0_0_0_10[7:0]  ), //o
    .io_outputs_7_payload_0_0_0_11    (streamDemux_2_io_outputs_7_payload_0_0_0_11[7:0]  ), //o
    .io_outputs_7_payload_0_0_0_12    (streamDemux_2_io_outputs_7_payload_0_0_0_12[7:0]  ), //o
    .io_outputs_7_payload_0_0_0_13    (streamDemux_2_io_outputs_7_payload_0_0_0_13[7:0]  ), //o
    .io_outputs_7_payload_0_0_0_14    (streamDemux_2_io_outputs_7_payload_0_0_0_14[7:0]  ), //o
    .io_outputs_7_payload_0_0_0_15    (streamDemux_2_io_outputs_7_payload_0_0_0_15[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_0     (streamDemux_2_io_outputs_7_payload_0_0_1_0[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_1     (streamDemux_2_io_outputs_7_payload_0_0_1_1[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_2     (streamDemux_2_io_outputs_7_payload_0_0_1_2[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_3     (streamDemux_2_io_outputs_7_payload_0_0_1_3[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_4     (streamDemux_2_io_outputs_7_payload_0_0_1_4[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_5     (streamDemux_2_io_outputs_7_payload_0_0_1_5[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_6     (streamDemux_2_io_outputs_7_payload_0_0_1_6[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_7     (streamDemux_2_io_outputs_7_payload_0_0_1_7[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_8     (streamDemux_2_io_outputs_7_payload_0_0_1_8[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_9     (streamDemux_2_io_outputs_7_payload_0_0_1_9[7:0]   ), //o
    .io_outputs_7_payload_0_0_1_10    (streamDemux_2_io_outputs_7_payload_0_0_1_10[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_11    (streamDemux_2_io_outputs_7_payload_0_0_1_11[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_12    (streamDemux_2_io_outputs_7_payload_0_0_1_12[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_13    (streamDemux_2_io_outputs_7_payload_0_0_1_13[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_14    (streamDemux_2_io_outputs_7_payload_0_0_1_14[7:0]  ), //o
    .io_outputs_7_payload_0_0_1_15    (streamDemux_2_io_outputs_7_payload_0_0_1_15[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_0     (streamDemux_2_io_outputs_7_payload_0_0_2_0[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_1     (streamDemux_2_io_outputs_7_payload_0_0_2_1[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_2     (streamDemux_2_io_outputs_7_payload_0_0_2_2[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_3     (streamDemux_2_io_outputs_7_payload_0_0_2_3[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_4     (streamDemux_2_io_outputs_7_payload_0_0_2_4[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_5     (streamDemux_2_io_outputs_7_payload_0_0_2_5[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_6     (streamDemux_2_io_outputs_7_payload_0_0_2_6[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_7     (streamDemux_2_io_outputs_7_payload_0_0_2_7[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_8     (streamDemux_2_io_outputs_7_payload_0_0_2_8[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_9     (streamDemux_2_io_outputs_7_payload_0_0_2_9[7:0]   ), //o
    .io_outputs_7_payload_0_0_2_10    (streamDemux_2_io_outputs_7_payload_0_0_2_10[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_11    (streamDemux_2_io_outputs_7_payload_0_0_2_11[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_12    (streamDemux_2_io_outputs_7_payload_0_0_2_12[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_13    (streamDemux_2_io_outputs_7_payload_0_0_2_13[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_14    (streamDemux_2_io_outputs_7_payload_0_0_2_14[7:0]  ), //o
    .io_outputs_7_payload_0_0_2_15    (streamDemux_2_io_outputs_7_payload_0_0_2_15[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_0     (streamDemux_2_io_outputs_7_payload_0_1_0_0[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_1     (streamDemux_2_io_outputs_7_payload_0_1_0_1[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_2     (streamDemux_2_io_outputs_7_payload_0_1_0_2[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_3     (streamDemux_2_io_outputs_7_payload_0_1_0_3[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_4     (streamDemux_2_io_outputs_7_payload_0_1_0_4[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_5     (streamDemux_2_io_outputs_7_payload_0_1_0_5[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_6     (streamDemux_2_io_outputs_7_payload_0_1_0_6[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_7     (streamDemux_2_io_outputs_7_payload_0_1_0_7[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_8     (streamDemux_2_io_outputs_7_payload_0_1_0_8[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_9     (streamDemux_2_io_outputs_7_payload_0_1_0_9[7:0]   ), //o
    .io_outputs_7_payload_0_1_0_10    (streamDemux_2_io_outputs_7_payload_0_1_0_10[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_11    (streamDemux_2_io_outputs_7_payload_0_1_0_11[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_12    (streamDemux_2_io_outputs_7_payload_0_1_0_12[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_13    (streamDemux_2_io_outputs_7_payload_0_1_0_13[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_14    (streamDemux_2_io_outputs_7_payload_0_1_0_14[7:0]  ), //o
    .io_outputs_7_payload_0_1_0_15    (streamDemux_2_io_outputs_7_payload_0_1_0_15[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_0     (streamDemux_2_io_outputs_7_payload_0_1_1_0[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_1     (streamDemux_2_io_outputs_7_payload_0_1_1_1[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_2     (streamDemux_2_io_outputs_7_payload_0_1_1_2[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_3     (streamDemux_2_io_outputs_7_payload_0_1_1_3[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_4     (streamDemux_2_io_outputs_7_payload_0_1_1_4[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_5     (streamDemux_2_io_outputs_7_payload_0_1_1_5[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_6     (streamDemux_2_io_outputs_7_payload_0_1_1_6[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_7     (streamDemux_2_io_outputs_7_payload_0_1_1_7[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_8     (streamDemux_2_io_outputs_7_payload_0_1_1_8[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_9     (streamDemux_2_io_outputs_7_payload_0_1_1_9[7:0]   ), //o
    .io_outputs_7_payload_0_1_1_10    (streamDemux_2_io_outputs_7_payload_0_1_1_10[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_11    (streamDemux_2_io_outputs_7_payload_0_1_1_11[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_12    (streamDemux_2_io_outputs_7_payload_0_1_1_12[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_13    (streamDemux_2_io_outputs_7_payload_0_1_1_13[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_14    (streamDemux_2_io_outputs_7_payload_0_1_1_14[7:0]  ), //o
    .io_outputs_7_payload_0_1_1_15    (streamDemux_2_io_outputs_7_payload_0_1_1_15[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_0     (streamDemux_2_io_outputs_7_payload_0_1_2_0[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_1     (streamDemux_2_io_outputs_7_payload_0_1_2_1[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_2     (streamDemux_2_io_outputs_7_payload_0_1_2_2[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_3     (streamDemux_2_io_outputs_7_payload_0_1_2_3[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_4     (streamDemux_2_io_outputs_7_payload_0_1_2_4[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_5     (streamDemux_2_io_outputs_7_payload_0_1_2_5[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_6     (streamDemux_2_io_outputs_7_payload_0_1_2_6[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_7     (streamDemux_2_io_outputs_7_payload_0_1_2_7[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_8     (streamDemux_2_io_outputs_7_payload_0_1_2_8[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_9     (streamDemux_2_io_outputs_7_payload_0_1_2_9[7:0]   ), //o
    .io_outputs_7_payload_0_1_2_10    (streamDemux_2_io_outputs_7_payload_0_1_2_10[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_11    (streamDemux_2_io_outputs_7_payload_0_1_2_11[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_12    (streamDemux_2_io_outputs_7_payload_0_1_2_12[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_13    (streamDemux_2_io_outputs_7_payload_0_1_2_13[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_14    (streamDemux_2_io_outputs_7_payload_0_1_2_14[7:0]  ), //o
    .io_outputs_7_payload_0_1_2_15    (streamDemux_2_io_outputs_7_payload_0_1_2_15[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_0     (streamDemux_2_io_outputs_7_payload_0_2_0_0[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_1     (streamDemux_2_io_outputs_7_payload_0_2_0_1[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_2     (streamDemux_2_io_outputs_7_payload_0_2_0_2[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_3     (streamDemux_2_io_outputs_7_payload_0_2_0_3[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_4     (streamDemux_2_io_outputs_7_payload_0_2_0_4[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_5     (streamDemux_2_io_outputs_7_payload_0_2_0_5[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_6     (streamDemux_2_io_outputs_7_payload_0_2_0_6[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_7     (streamDemux_2_io_outputs_7_payload_0_2_0_7[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_8     (streamDemux_2_io_outputs_7_payload_0_2_0_8[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_9     (streamDemux_2_io_outputs_7_payload_0_2_0_9[7:0]   ), //o
    .io_outputs_7_payload_0_2_0_10    (streamDemux_2_io_outputs_7_payload_0_2_0_10[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_11    (streamDemux_2_io_outputs_7_payload_0_2_0_11[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_12    (streamDemux_2_io_outputs_7_payload_0_2_0_12[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_13    (streamDemux_2_io_outputs_7_payload_0_2_0_13[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_14    (streamDemux_2_io_outputs_7_payload_0_2_0_14[7:0]  ), //o
    .io_outputs_7_payload_0_2_0_15    (streamDemux_2_io_outputs_7_payload_0_2_0_15[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_0     (streamDemux_2_io_outputs_7_payload_0_2_1_0[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_1     (streamDemux_2_io_outputs_7_payload_0_2_1_1[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_2     (streamDemux_2_io_outputs_7_payload_0_2_1_2[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_3     (streamDemux_2_io_outputs_7_payload_0_2_1_3[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_4     (streamDemux_2_io_outputs_7_payload_0_2_1_4[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_5     (streamDemux_2_io_outputs_7_payload_0_2_1_5[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_6     (streamDemux_2_io_outputs_7_payload_0_2_1_6[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_7     (streamDemux_2_io_outputs_7_payload_0_2_1_7[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_8     (streamDemux_2_io_outputs_7_payload_0_2_1_8[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_9     (streamDemux_2_io_outputs_7_payload_0_2_1_9[7:0]   ), //o
    .io_outputs_7_payload_0_2_1_10    (streamDemux_2_io_outputs_7_payload_0_2_1_10[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_11    (streamDemux_2_io_outputs_7_payload_0_2_1_11[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_12    (streamDemux_2_io_outputs_7_payload_0_2_1_12[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_13    (streamDemux_2_io_outputs_7_payload_0_2_1_13[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_14    (streamDemux_2_io_outputs_7_payload_0_2_1_14[7:0]  ), //o
    .io_outputs_7_payload_0_2_1_15    (streamDemux_2_io_outputs_7_payload_0_2_1_15[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_0     (streamDemux_2_io_outputs_7_payload_0_2_2_0[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_1     (streamDemux_2_io_outputs_7_payload_0_2_2_1[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_2     (streamDemux_2_io_outputs_7_payload_0_2_2_2[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_3     (streamDemux_2_io_outputs_7_payload_0_2_2_3[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_4     (streamDemux_2_io_outputs_7_payload_0_2_2_4[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_5     (streamDemux_2_io_outputs_7_payload_0_2_2_5[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_6     (streamDemux_2_io_outputs_7_payload_0_2_2_6[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_7     (streamDemux_2_io_outputs_7_payload_0_2_2_7[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_8     (streamDemux_2_io_outputs_7_payload_0_2_2_8[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_9     (streamDemux_2_io_outputs_7_payload_0_2_2_9[7:0]   ), //o
    .io_outputs_7_payload_0_2_2_10    (streamDemux_2_io_outputs_7_payload_0_2_2_10[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_11    (streamDemux_2_io_outputs_7_payload_0_2_2_11[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_12    (streamDemux_2_io_outputs_7_payload_0_2_2_12[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_13    (streamDemux_2_io_outputs_7_payload_0_2_2_13[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_14    (streamDemux_2_io_outputs_7_payload_0_2_2_14[7:0]  ), //o
    .io_outputs_7_payload_0_2_2_15    (streamDemux_2_io_outputs_7_payload_0_2_2_15[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_0     (streamDemux_2_io_outputs_7_payload_1_0_0_0[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_1     (streamDemux_2_io_outputs_7_payload_1_0_0_1[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_2     (streamDemux_2_io_outputs_7_payload_1_0_0_2[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_3     (streamDemux_2_io_outputs_7_payload_1_0_0_3[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_4     (streamDemux_2_io_outputs_7_payload_1_0_0_4[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_5     (streamDemux_2_io_outputs_7_payload_1_0_0_5[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_6     (streamDemux_2_io_outputs_7_payload_1_0_0_6[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_7     (streamDemux_2_io_outputs_7_payload_1_0_0_7[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_8     (streamDemux_2_io_outputs_7_payload_1_0_0_8[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_9     (streamDemux_2_io_outputs_7_payload_1_0_0_9[7:0]   ), //o
    .io_outputs_7_payload_1_0_0_10    (streamDemux_2_io_outputs_7_payload_1_0_0_10[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_11    (streamDemux_2_io_outputs_7_payload_1_0_0_11[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_12    (streamDemux_2_io_outputs_7_payload_1_0_0_12[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_13    (streamDemux_2_io_outputs_7_payload_1_0_0_13[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_14    (streamDemux_2_io_outputs_7_payload_1_0_0_14[7:0]  ), //o
    .io_outputs_7_payload_1_0_0_15    (streamDemux_2_io_outputs_7_payload_1_0_0_15[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_0     (streamDemux_2_io_outputs_7_payload_1_0_1_0[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_1     (streamDemux_2_io_outputs_7_payload_1_0_1_1[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_2     (streamDemux_2_io_outputs_7_payload_1_0_1_2[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_3     (streamDemux_2_io_outputs_7_payload_1_0_1_3[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_4     (streamDemux_2_io_outputs_7_payload_1_0_1_4[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_5     (streamDemux_2_io_outputs_7_payload_1_0_1_5[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_6     (streamDemux_2_io_outputs_7_payload_1_0_1_6[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_7     (streamDemux_2_io_outputs_7_payload_1_0_1_7[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_8     (streamDemux_2_io_outputs_7_payload_1_0_1_8[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_9     (streamDemux_2_io_outputs_7_payload_1_0_1_9[7:0]   ), //o
    .io_outputs_7_payload_1_0_1_10    (streamDemux_2_io_outputs_7_payload_1_0_1_10[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_11    (streamDemux_2_io_outputs_7_payload_1_0_1_11[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_12    (streamDemux_2_io_outputs_7_payload_1_0_1_12[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_13    (streamDemux_2_io_outputs_7_payload_1_0_1_13[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_14    (streamDemux_2_io_outputs_7_payload_1_0_1_14[7:0]  ), //o
    .io_outputs_7_payload_1_0_1_15    (streamDemux_2_io_outputs_7_payload_1_0_1_15[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_0     (streamDemux_2_io_outputs_7_payload_1_0_2_0[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_1     (streamDemux_2_io_outputs_7_payload_1_0_2_1[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_2     (streamDemux_2_io_outputs_7_payload_1_0_2_2[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_3     (streamDemux_2_io_outputs_7_payload_1_0_2_3[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_4     (streamDemux_2_io_outputs_7_payload_1_0_2_4[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_5     (streamDemux_2_io_outputs_7_payload_1_0_2_5[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_6     (streamDemux_2_io_outputs_7_payload_1_0_2_6[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_7     (streamDemux_2_io_outputs_7_payload_1_0_2_7[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_8     (streamDemux_2_io_outputs_7_payload_1_0_2_8[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_9     (streamDemux_2_io_outputs_7_payload_1_0_2_9[7:0]   ), //o
    .io_outputs_7_payload_1_0_2_10    (streamDemux_2_io_outputs_7_payload_1_0_2_10[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_11    (streamDemux_2_io_outputs_7_payload_1_0_2_11[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_12    (streamDemux_2_io_outputs_7_payload_1_0_2_12[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_13    (streamDemux_2_io_outputs_7_payload_1_0_2_13[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_14    (streamDemux_2_io_outputs_7_payload_1_0_2_14[7:0]  ), //o
    .io_outputs_7_payload_1_0_2_15    (streamDemux_2_io_outputs_7_payload_1_0_2_15[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_0     (streamDemux_2_io_outputs_7_payload_1_1_0_0[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_1     (streamDemux_2_io_outputs_7_payload_1_1_0_1[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_2     (streamDemux_2_io_outputs_7_payload_1_1_0_2[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_3     (streamDemux_2_io_outputs_7_payload_1_1_0_3[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_4     (streamDemux_2_io_outputs_7_payload_1_1_0_4[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_5     (streamDemux_2_io_outputs_7_payload_1_1_0_5[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_6     (streamDemux_2_io_outputs_7_payload_1_1_0_6[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_7     (streamDemux_2_io_outputs_7_payload_1_1_0_7[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_8     (streamDemux_2_io_outputs_7_payload_1_1_0_8[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_9     (streamDemux_2_io_outputs_7_payload_1_1_0_9[7:0]   ), //o
    .io_outputs_7_payload_1_1_0_10    (streamDemux_2_io_outputs_7_payload_1_1_0_10[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_11    (streamDemux_2_io_outputs_7_payload_1_1_0_11[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_12    (streamDemux_2_io_outputs_7_payload_1_1_0_12[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_13    (streamDemux_2_io_outputs_7_payload_1_1_0_13[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_14    (streamDemux_2_io_outputs_7_payload_1_1_0_14[7:0]  ), //o
    .io_outputs_7_payload_1_1_0_15    (streamDemux_2_io_outputs_7_payload_1_1_0_15[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_0     (streamDemux_2_io_outputs_7_payload_1_1_1_0[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_1     (streamDemux_2_io_outputs_7_payload_1_1_1_1[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_2     (streamDemux_2_io_outputs_7_payload_1_1_1_2[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_3     (streamDemux_2_io_outputs_7_payload_1_1_1_3[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_4     (streamDemux_2_io_outputs_7_payload_1_1_1_4[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_5     (streamDemux_2_io_outputs_7_payload_1_1_1_5[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_6     (streamDemux_2_io_outputs_7_payload_1_1_1_6[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_7     (streamDemux_2_io_outputs_7_payload_1_1_1_7[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_8     (streamDemux_2_io_outputs_7_payload_1_1_1_8[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_9     (streamDemux_2_io_outputs_7_payload_1_1_1_9[7:0]   ), //o
    .io_outputs_7_payload_1_1_1_10    (streamDemux_2_io_outputs_7_payload_1_1_1_10[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_11    (streamDemux_2_io_outputs_7_payload_1_1_1_11[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_12    (streamDemux_2_io_outputs_7_payload_1_1_1_12[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_13    (streamDemux_2_io_outputs_7_payload_1_1_1_13[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_14    (streamDemux_2_io_outputs_7_payload_1_1_1_14[7:0]  ), //o
    .io_outputs_7_payload_1_1_1_15    (streamDemux_2_io_outputs_7_payload_1_1_1_15[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_0     (streamDemux_2_io_outputs_7_payload_1_1_2_0[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_1     (streamDemux_2_io_outputs_7_payload_1_1_2_1[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_2     (streamDemux_2_io_outputs_7_payload_1_1_2_2[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_3     (streamDemux_2_io_outputs_7_payload_1_1_2_3[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_4     (streamDemux_2_io_outputs_7_payload_1_1_2_4[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_5     (streamDemux_2_io_outputs_7_payload_1_1_2_5[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_6     (streamDemux_2_io_outputs_7_payload_1_1_2_6[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_7     (streamDemux_2_io_outputs_7_payload_1_1_2_7[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_8     (streamDemux_2_io_outputs_7_payload_1_1_2_8[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_9     (streamDemux_2_io_outputs_7_payload_1_1_2_9[7:0]   ), //o
    .io_outputs_7_payload_1_1_2_10    (streamDemux_2_io_outputs_7_payload_1_1_2_10[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_11    (streamDemux_2_io_outputs_7_payload_1_1_2_11[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_12    (streamDemux_2_io_outputs_7_payload_1_1_2_12[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_13    (streamDemux_2_io_outputs_7_payload_1_1_2_13[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_14    (streamDemux_2_io_outputs_7_payload_1_1_2_14[7:0]  ), //o
    .io_outputs_7_payload_1_1_2_15    (streamDemux_2_io_outputs_7_payload_1_1_2_15[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_0     (streamDemux_2_io_outputs_7_payload_1_2_0_0[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_1     (streamDemux_2_io_outputs_7_payload_1_2_0_1[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_2     (streamDemux_2_io_outputs_7_payload_1_2_0_2[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_3     (streamDemux_2_io_outputs_7_payload_1_2_0_3[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_4     (streamDemux_2_io_outputs_7_payload_1_2_0_4[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_5     (streamDemux_2_io_outputs_7_payload_1_2_0_5[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_6     (streamDemux_2_io_outputs_7_payload_1_2_0_6[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_7     (streamDemux_2_io_outputs_7_payload_1_2_0_7[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_8     (streamDemux_2_io_outputs_7_payload_1_2_0_8[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_9     (streamDemux_2_io_outputs_7_payload_1_2_0_9[7:0]   ), //o
    .io_outputs_7_payload_1_2_0_10    (streamDemux_2_io_outputs_7_payload_1_2_0_10[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_11    (streamDemux_2_io_outputs_7_payload_1_2_0_11[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_12    (streamDemux_2_io_outputs_7_payload_1_2_0_12[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_13    (streamDemux_2_io_outputs_7_payload_1_2_0_13[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_14    (streamDemux_2_io_outputs_7_payload_1_2_0_14[7:0]  ), //o
    .io_outputs_7_payload_1_2_0_15    (streamDemux_2_io_outputs_7_payload_1_2_0_15[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_0     (streamDemux_2_io_outputs_7_payload_1_2_1_0[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_1     (streamDemux_2_io_outputs_7_payload_1_2_1_1[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_2     (streamDemux_2_io_outputs_7_payload_1_2_1_2[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_3     (streamDemux_2_io_outputs_7_payload_1_2_1_3[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_4     (streamDemux_2_io_outputs_7_payload_1_2_1_4[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_5     (streamDemux_2_io_outputs_7_payload_1_2_1_5[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_6     (streamDemux_2_io_outputs_7_payload_1_2_1_6[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_7     (streamDemux_2_io_outputs_7_payload_1_2_1_7[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_8     (streamDemux_2_io_outputs_7_payload_1_2_1_8[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_9     (streamDemux_2_io_outputs_7_payload_1_2_1_9[7:0]   ), //o
    .io_outputs_7_payload_1_2_1_10    (streamDemux_2_io_outputs_7_payload_1_2_1_10[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_11    (streamDemux_2_io_outputs_7_payload_1_2_1_11[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_12    (streamDemux_2_io_outputs_7_payload_1_2_1_12[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_13    (streamDemux_2_io_outputs_7_payload_1_2_1_13[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_14    (streamDemux_2_io_outputs_7_payload_1_2_1_14[7:0]  ), //o
    .io_outputs_7_payload_1_2_1_15    (streamDemux_2_io_outputs_7_payload_1_2_1_15[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_0     (streamDemux_2_io_outputs_7_payload_1_2_2_0[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_1     (streamDemux_2_io_outputs_7_payload_1_2_2_1[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_2     (streamDemux_2_io_outputs_7_payload_1_2_2_2[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_3     (streamDemux_2_io_outputs_7_payload_1_2_2_3[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_4     (streamDemux_2_io_outputs_7_payload_1_2_2_4[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_5     (streamDemux_2_io_outputs_7_payload_1_2_2_5[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_6     (streamDemux_2_io_outputs_7_payload_1_2_2_6[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_7     (streamDemux_2_io_outputs_7_payload_1_2_2_7[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_8     (streamDemux_2_io_outputs_7_payload_1_2_2_8[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_9     (streamDemux_2_io_outputs_7_payload_1_2_2_9[7:0]   ), //o
    .io_outputs_7_payload_1_2_2_10    (streamDemux_2_io_outputs_7_payload_1_2_2_10[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_11    (streamDemux_2_io_outputs_7_payload_1_2_2_11[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_12    (streamDemux_2_io_outputs_7_payload_1_2_2_12[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_13    (streamDemux_2_io_outputs_7_payload_1_2_2_13[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_14    (streamDemux_2_io_outputs_7_payload_1_2_2_14[7:0]  ), //o
    .io_outputs_7_payload_1_2_2_15    (streamDemux_2_io_outputs_7_payload_1_2_2_15[7:0]  )  //o
  );
  EventM2sPipes_8 eventM2sPipes_9 (
    .eventIn_valid     (accOutputsJoin_valid            ), //i
    .eventIn_ready     (eventM2sPipes_9_eventIn_ready   ), //o
    .eventOut_valid    (eventM2sPipes_9_eventOut_valid  ), //o
    .eventOut_ready    (postProcessOutputs_ready        ), //i
    .CEs_0             (eventM2sPipes_9_CEs_0           ), //o
    .CEs_1             (eventM2sPipes_9_CEs_1           ), //o
    .CEs_2             (eventM2sPipes_9_CEs_2           ), //o
    .CEs_3             (eventM2sPipes_9_CEs_3           ), //o
    .CEs_4             (eventM2sPipes_9_CEs_4           ), //o
    .CEs_5             (eventM2sPipes_9_CEs_5           ), //o
    .clk               (clk                             ), //i
    .reset             (reset                           )  //i
  );
  ScalerINT16 scalerINT16_16 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_0[23:0]  ), //i
    .dout          (scalerINT16_16_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_17 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_1[23:0]  ), //i
    .dout          (scalerINT16_17_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_18 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_2[23:0]  ), //i
    .dout          (scalerINT16_18_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_19 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_3[23:0]  ), //i
    .dout          (scalerINT16_19_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_20 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_4[23:0]  ), //i
    .dout          (scalerINT16_20_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_21 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_5[23:0]  ), //i
    .dout          (scalerINT16_21_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_22 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_6[23:0]  ), //i
    .dout          (scalerINT16_22_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_23 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_7[23:0]  ), //i
    .dout          (scalerINT16_23_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_24 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_8[23:0]  ), //i
    .dout          (scalerINT16_24_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_25 (
    .scalerBase    (scaleBase[15:0]                                  ), //i
    .scalerExpr    (scaleExpr[5:0]                                   ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                            ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                            ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                            ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                            ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                            ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                            ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_9[23:0]  ), //i
    .dout          (scalerINT16_25_dout[7:0]                         ), //o
    .clk           (clk                                              ), //i
    .reset         (reset                                            )  //i
  );
  ScalerINT16 scalerINT16_26 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_10[23:0]  ), //i
    .dout          (scalerINT16_26_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  ScalerINT16 scalerINT16_27 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_11[23:0]  ), //i
    .dout          (scalerINT16_27_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  ScalerINT16 scalerINT16_28 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_12[23:0]  ), //i
    .dout          (scalerINT16_28_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  ScalerINT16 scalerINT16_29 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_13[23:0]  ), //i
    .dout          (scalerINT16_29_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  ScalerINT16 scalerINT16_30 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_14[23:0]  ), //i
    .dout          (scalerINT16_30_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  ScalerINT16 scalerINT16_31 (
    .scalerBase    (scaleBase[15:0]                                   ), //i
    .scalerExpr    (scaleExpr[5:0]                                    ), //i
    .CEs_0         (eventM2sPipes_9_CEs_0                             ), //i
    .CEs_1         (eventM2sPipes_9_CEs_1                             ), //i
    .CEs_2         (eventM2sPipes_9_CEs_2                             ), //i
    .CEs_3         (eventM2sPipes_9_CEs_3                             ), //i
    .CEs_4         (eventM2sPipes_9_CEs_4                             ), //i
    .CEs_5         (eventM2sPipes_9_CEs_5                             ), //i
    .din           (accOutputsJoin_payload_frame_line_pixel_15[23:0]  ), //i
    .dout          (scalerINT16_31_dout[7:0]                          ), //o
    .clk           (clk                                               ), //i
    .reset         (reset                                             )  //i
  );
  StreamDemux_1 streamDemux_3 (
    .io_select                                    (streamDemux_3_io_select                                      ), //i
    .io_input_valid                               (postProcessOutputs_valid                                     ), //i
    .io_input_ready                               (streamDemux_3_io_input_ready                                 ), //o
    .io_input_payload_frame_line_pixel_0          (postProcessOutputs_payload_frame_line_pixel_0[7:0]           ), //i
    .io_input_payload_frame_line_pixel_1          (postProcessOutputs_payload_frame_line_pixel_1[7:0]           ), //i
    .io_input_payload_frame_line_pixel_2          (postProcessOutputs_payload_frame_line_pixel_2[7:0]           ), //i
    .io_input_payload_frame_line_pixel_3          (postProcessOutputs_payload_frame_line_pixel_3[7:0]           ), //i
    .io_input_payload_frame_line_pixel_4          (postProcessOutputs_payload_frame_line_pixel_4[7:0]           ), //i
    .io_input_payload_frame_line_pixel_5          (postProcessOutputs_payload_frame_line_pixel_5[7:0]           ), //i
    .io_input_payload_frame_line_pixel_6          (postProcessOutputs_payload_frame_line_pixel_6[7:0]           ), //i
    .io_input_payload_frame_line_pixel_7          (postProcessOutputs_payload_frame_line_pixel_7[7:0]           ), //i
    .io_input_payload_frame_line_pixel_8          (postProcessOutputs_payload_frame_line_pixel_8[7:0]           ), //i
    .io_input_payload_frame_line_pixel_9          (postProcessOutputs_payload_frame_line_pixel_9[7:0]           ), //i
    .io_input_payload_frame_line_pixel_10         (postProcessOutputs_payload_frame_line_pixel_10[7:0]          ), //i
    .io_input_payload_frame_line_pixel_11         (postProcessOutputs_payload_frame_line_pixel_11[7:0]          ), //i
    .io_input_payload_frame_line_pixel_12         (postProcessOutputs_payload_frame_line_pixel_12[7:0]          ), //i
    .io_input_payload_frame_line_pixel_13         (postProcessOutputs_payload_frame_line_pixel_13[7:0]          ), //i
    .io_input_payload_frame_line_pixel_14         (postProcessOutputs_payload_frame_line_pixel_14[7:0]          ), //i
    .io_input_payload_frame_line_pixel_15         (postProcessOutputs_payload_frame_line_pixel_15[7:0]          ), //i
    .io_input_payload_frame_line_endOfLine        (postProcessOutputs_payload_frame_line_endOfLine              ), //i
    .io_input_payload_frame_endOfFrame            (postProcessOutputs_payload_frame_endOfFrame                  ), //i
    .io_input_payload_endOfPack                   (postProcessOutputs_payload_endOfPack                         ), //i
    .io_outputs_0_valid                           (streamDemux_3_io_outputs_0_valid                             ), //o
    .io_outputs_0_ready                           (streamMux_1_io_inputs_0_ready                                ), //i
    .io_outputs_0_payload_frame_line_pixel_0      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_3      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_4      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_5      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_6      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_7      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_8      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_9      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_10     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_11     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_12     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_13     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_14     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_15     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_endOfLine    (streamDemux_3_io_outputs_0_payload_frame_line_endOfLine      ), //o
    .io_outputs_0_payload_frame_endOfFrame        (streamDemux_3_io_outputs_0_payload_frame_endOfFrame          ), //o
    .io_outputs_0_payload_endOfPack               (streamDemux_3_io_outputs_0_payload_endOfPack                 ), //o
    .io_outputs_1_valid                           (streamDemux_3_io_outputs_1_valid                             ), //o
    .io_outputs_1_ready                           (pool_videoIn_ready                                           ), //i
    .io_outputs_1_payload_frame_line_pixel_0      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_3      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_4      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_5      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_6      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_7      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_8      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_9      (streamDemux_3_io_outputs_1_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_10     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_11     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_12     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_13     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_14     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_15     (streamDemux_3_io_outputs_1_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_endOfLine    (streamDemux_3_io_outputs_1_payload_frame_line_endOfLine      ), //o
    .io_outputs_1_payload_frame_endOfFrame        (streamDemux_3_io_outputs_1_payload_frame_endOfFrame          ), //o
    .io_outputs_1_payload_endOfPack               (streamDemux_3_io_outputs_1_payload_endOfPack                 )  //o
  );
  StreamMux streamMux_1 (
    .io_select                                   (streamMux_1_io_select                                        ), //i
    .io_inputs_0_valid                           (streamDemux_3_io_outputs_0_valid                             ), //i
    .io_inputs_0_ready                           (streamMux_1_io_inputs_0_ready                                ), //o
    .io_inputs_0_payload_frame_line_pixel_0      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_0[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_1      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_1[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_2      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_2[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_3      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_3[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_4      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_4[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_5      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_5[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_6      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_6[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_7      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_7[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_8      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_8[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_9      (streamDemux_3_io_outputs_0_payload_frame_line_pixel_9[7:0]   ), //i
    .io_inputs_0_payload_frame_line_pixel_10     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_10[7:0]  ), //i
    .io_inputs_0_payload_frame_line_pixel_11     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_11[7:0]  ), //i
    .io_inputs_0_payload_frame_line_pixel_12     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_12[7:0]  ), //i
    .io_inputs_0_payload_frame_line_pixel_13     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_13[7:0]  ), //i
    .io_inputs_0_payload_frame_line_pixel_14     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_14[7:0]  ), //i
    .io_inputs_0_payload_frame_line_pixel_15     (streamDemux_3_io_outputs_0_payload_frame_line_pixel_15[7:0]  ), //i
    .io_inputs_0_payload_frame_line_endOfLine    (streamDemux_3_io_outputs_0_payload_frame_line_endOfLine      ), //i
    .io_inputs_0_payload_frame_endOfFrame        (streamDemux_3_io_outputs_0_payload_frame_endOfFrame          ), //i
    .io_inputs_0_payload_endOfPack               (streamDemux_3_io_outputs_0_payload_endOfPack                 ), //i
    .io_inputs_1_valid                           (pool_videoOut_valid                                          ), //i
    .io_inputs_1_ready                           (streamMux_1_io_inputs_1_ready                                ), //o
    .io_inputs_1_payload_frame_line_pixel_0      (pool_videoOut_payload_frame_line_pixel_0[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_1      (pool_videoOut_payload_frame_line_pixel_1[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_2      (pool_videoOut_payload_frame_line_pixel_2[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_3      (pool_videoOut_payload_frame_line_pixel_3[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_4      (pool_videoOut_payload_frame_line_pixel_4[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_5      (pool_videoOut_payload_frame_line_pixel_5[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_6      (pool_videoOut_payload_frame_line_pixel_6[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_7      (pool_videoOut_payload_frame_line_pixel_7[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_8      (pool_videoOut_payload_frame_line_pixel_8[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_9      (pool_videoOut_payload_frame_line_pixel_9[7:0]                ), //i
    .io_inputs_1_payload_frame_line_pixel_10     (pool_videoOut_payload_frame_line_pixel_10[7:0]               ), //i
    .io_inputs_1_payload_frame_line_pixel_11     (pool_videoOut_payload_frame_line_pixel_11[7:0]               ), //i
    .io_inputs_1_payload_frame_line_pixel_12     (pool_videoOut_payload_frame_line_pixel_12[7:0]               ), //i
    .io_inputs_1_payload_frame_line_pixel_13     (pool_videoOut_payload_frame_line_pixel_13[7:0]               ), //i
    .io_inputs_1_payload_frame_line_pixel_14     (pool_videoOut_payload_frame_line_pixel_14[7:0]               ), //i
    .io_inputs_1_payload_frame_line_pixel_15     (pool_videoOut_payload_frame_line_pixel_15[7:0]               ), //i
    .io_inputs_1_payload_frame_line_endOfLine    (pool_videoOut_payload_frame_line_endOfLine                   ), //i
    .io_inputs_1_payload_frame_endOfFrame        (pool_videoOut_payload_frame_endOfFrame                       ), //i
    .io_inputs_1_payload_endOfPack               (pool_videoOut_payload_endOfPack                              ), //i
    .io_output_valid                             (streamMux_1_io_output_valid                                  ), //o
    .io_output_ready                             (streamMux_1_io_output_translated_ready                       ), //i
    .io_output_payload_frame_line_pixel_0        (streamMux_1_io_output_payload_frame_line_pixel_0[7:0]        ), //o
    .io_output_payload_frame_line_pixel_1        (streamMux_1_io_output_payload_frame_line_pixel_1[7:0]        ), //o
    .io_output_payload_frame_line_pixel_2        (streamMux_1_io_output_payload_frame_line_pixel_2[7:0]        ), //o
    .io_output_payload_frame_line_pixel_3        (streamMux_1_io_output_payload_frame_line_pixel_3[7:0]        ), //o
    .io_output_payload_frame_line_pixel_4        (streamMux_1_io_output_payload_frame_line_pixel_4[7:0]        ), //o
    .io_output_payload_frame_line_pixel_5        (streamMux_1_io_output_payload_frame_line_pixel_5[7:0]        ), //o
    .io_output_payload_frame_line_pixel_6        (streamMux_1_io_output_payload_frame_line_pixel_6[7:0]        ), //o
    .io_output_payload_frame_line_pixel_7        (streamMux_1_io_output_payload_frame_line_pixel_7[7:0]        ), //o
    .io_output_payload_frame_line_pixel_8        (streamMux_1_io_output_payload_frame_line_pixel_8[7:0]        ), //o
    .io_output_payload_frame_line_pixel_9        (streamMux_1_io_output_payload_frame_line_pixel_9[7:0]        ), //o
    .io_output_payload_frame_line_pixel_10       (streamMux_1_io_output_payload_frame_line_pixel_10[7:0]       ), //o
    .io_output_payload_frame_line_pixel_11       (streamMux_1_io_output_payload_frame_line_pixel_11[7:0]       ), //o
    .io_output_payload_frame_line_pixel_12       (streamMux_1_io_output_payload_frame_line_pixel_12[7:0]       ), //o
    .io_output_payload_frame_line_pixel_13       (streamMux_1_io_output_payload_frame_line_pixel_13[7:0]       ), //o
    .io_output_payload_frame_line_pixel_14       (streamMux_1_io_output_payload_frame_line_pixel_14[7:0]       ), //o
    .io_output_payload_frame_line_pixel_15       (streamMux_1_io_output_payload_frame_line_pixel_15[7:0]       ), //o
    .io_output_payload_frame_line_endOfLine      (streamMux_1_io_output_payload_frame_line_endOfLine           ), //o
    .io_output_payload_frame_endOfFrame          (streamMux_1_io_output_payload_frame_endOfFrame               ), //o
    .io_output_payload_endOfPack                 (streamMux_1_io_output_payload_endOfPack                      )  //o
  );
  always @(*) begin
    case(tmp_funcTable_ready_2)
      4'b0000 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[7 : 0];
      4'b0001 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[15 : 8];
      4'b0010 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[23 : 16];
      4'b0011 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[31 : 24];
      4'b0100 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[39 : 32];
      4'b0101 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[47 : 40];
      4'b0110 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[55 : 48];
      4'b0111 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[63 : 56];
      4'b1000 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[71 : 64];
      4'b1001 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[79 : 72];
      4'b1010 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[87 : 80];
      4'b1011 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[95 : 88];
      4'b1100 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[103 : 96];
      4'b1101 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[111 : 104];
      4'b1110 : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[119 : 112];
      default : tmp_tableAdapted_payload_1 = tmp_tableAdapted_payload[127 : 120];
    endcase
  end

  assign inputChannelSpilt_valid = inputs_valid;
  assign inputs_ready = inputChannelSpilt_ready;
  assign tmp_inputChannelSpilt_payload_0 = inputs_payload;
  assign inputChannelSpilt_payload_0 = tmp_inputChannelSpilt_payload_0[7 : 0];
  assign inputChannelSpilt_payload_1 = tmp_inputChannelSpilt_payload_0[15 : 8];
  assign inputChannelSpilt_payload_2 = tmp_inputChannelSpilt_payload_0[23 : 16];
  assign inputChannelSpilt_payload_3 = tmp_inputChannelSpilt_payload_0[31 : 24];
  assign inputChannelSpilt_payload_4 = tmp_inputChannelSpilt_payload_0[39 : 32];
  assign inputChannelSpilt_payload_5 = tmp_inputChannelSpilt_payload_0[47 : 40];
  assign inputChannelSpilt_payload_6 = tmp_inputChannelSpilt_payload_0[55 : 48];
  assign inputChannelSpilt_payload_7 = tmp_inputChannelSpilt_payload_0[63 : 56];
  assign inputChannelSpilt_payload_8 = tmp_inputChannelSpilt_payload_0[71 : 64];
  assign inputChannelSpilt_payload_9 = tmp_inputChannelSpilt_payload_0[79 : 72];
  assign inputChannelSpilt_payload_10 = tmp_inputChannelSpilt_payload_0[87 : 80];
  assign inputChannelSpilt_payload_11 = tmp_inputChannelSpilt_payload_0[95 : 88];
  assign inputChannelSpilt_payload_12 = tmp_inputChannelSpilt_payload_0[103 : 96];
  assign inputChannelSpilt_payload_13 = tmp_inputChannelSpilt_payload_0[111 : 104];
  assign inputChannelSpilt_payload_14 = tmp_inputChannelSpilt_payload_0[119 : 112];
  assign inputChannelSpilt_payload_15 = tmp_inputChannelSpilt_payload_0[127 : 120];
  assign inputChannelSpilt_translated_valid = inputChannelSpilt_valid;
  assign inputChannelSpilt_ready = inputChannelSpilt_translated_ready;
  assign inputChannelSpilt_translated_payload_0 = ($signed(inputChannelSpilt_payload_0) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_1 = ($signed(inputChannelSpilt_payload_1) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_2 = ($signed(inputChannelSpilt_payload_2) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_3 = ($signed(inputChannelSpilt_payload_3) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_4 = ($signed(inputChannelSpilt_payload_4) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_5 = ($signed(inputChannelSpilt_payload_5) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_6 = ($signed(inputChannelSpilt_payload_6) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_7 = ($signed(inputChannelSpilt_payload_7) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_8 = ($signed(inputChannelSpilt_payload_8) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_9 = ($signed(inputChannelSpilt_payload_9) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_10 = ($signed(inputChannelSpilt_payload_10) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_11 = ($signed(inputChannelSpilt_payload_11) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_12 = ($signed(inputChannelSpilt_payload_12) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_13 = ($signed(inputChannelSpilt_payload_13) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_14 = ($signed(inputChannelSpilt_payload_14) - $signed(inputZeroPoint));
  assign inputChannelSpilt_translated_payload_15 = ($signed(inputChannelSpilt_payload_15) - $signed(inputZeroPoint));
  always @(*) begin
    inputChannelSpilt_translated_ready = inputChannelSpilt_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      inputChannelSpilt_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! inputChannelSpilt_translated_m2sPipe_valid);
  assign inputChannelSpilt_translated_m2sPipe_valid = inputChannelSpilt_translated_rValid;
  assign inputChannelSpilt_translated_m2sPipe_payload_0 = inputChannelSpilt_translated_rData_0;
  assign inputChannelSpilt_translated_m2sPipe_payload_1 = inputChannelSpilt_translated_rData_1;
  assign inputChannelSpilt_translated_m2sPipe_payload_2 = inputChannelSpilt_translated_rData_2;
  assign inputChannelSpilt_translated_m2sPipe_payload_3 = inputChannelSpilt_translated_rData_3;
  assign inputChannelSpilt_translated_m2sPipe_payload_4 = inputChannelSpilt_translated_rData_4;
  assign inputChannelSpilt_translated_m2sPipe_payload_5 = inputChannelSpilt_translated_rData_5;
  assign inputChannelSpilt_translated_m2sPipe_payload_6 = inputChannelSpilt_translated_rData_6;
  assign inputChannelSpilt_translated_m2sPipe_payload_7 = inputChannelSpilt_translated_rData_7;
  assign inputChannelSpilt_translated_m2sPipe_payload_8 = inputChannelSpilt_translated_rData_8;
  assign inputChannelSpilt_translated_m2sPipe_payload_9 = inputChannelSpilt_translated_rData_9;
  assign inputChannelSpilt_translated_m2sPipe_payload_10 = inputChannelSpilt_translated_rData_10;
  assign inputChannelSpilt_translated_m2sPipe_payload_11 = inputChannelSpilt_translated_rData_11;
  assign inputChannelSpilt_translated_m2sPipe_payload_12 = inputChannelSpilt_translated_rData_12;
  assign inputChannelSpilt_translated_m2sPipe_payload_13 = inputChannelSpilt_translated_rData_13;
  assign inputChannelSpilt_translated_m2sPipe_payload_14 = inputChannelSpilt_translated_rData_14;
  assign inputChannelSpilt_translated_m2sPipe_payload_15 = inputChannelSpilt_translated_rData_15;
  assign inputChannelSpilt_translated_m2sPipe_fire = (inputChannelSpilt_translated_m2sPipe_valid && inputChannelSpilt_translated_m2sPipe_ready);
  always @(*) begin
    tmp_when_Utils_l503_2 = 1'b0;
    if(inputChannelSpilt_translated_m2sPipe_fire) begin
      tmp_when_Utils_l503_2 = 1'b1;
    end
  end

  always @(*) begin
    tmp_when_Utils_l503_3 = (tmp_when_Utils_l503_4 + tmp_tmp_when_Utils_l503_3);
    if(1'b0) begin
      tmp_when_Utils_l503_3 = 9'h0;
    end
  end

  assign when_Utils_l503 = (inputChannelSpilt_translated_m2sPipe_fire && tmp_when_Utils_l503);
  always @(*) begin
    tmp_when_Utils_l503_5 = 1'b0;
    if(when_Utils_l503) begin
      tmp_when_Utils_l503_5 = 1'b1;
    end
  end

  always @(*) begin
    tmp_when_Utils_l503_6 = (tmp_when_Utils_l503_7 + tmp_tmp_when_Utils_l503_6);
    if(1'b0) begin
      tmp_when_Utils_l503_6 = 9'h0;
    end
  end

  assign when_Utils_l503_1 = (inputChannelSpilt_translated_m2sPipe_fire && tmp_when_Utils_l503_1);
  always @(*) begin
    tmp_inputVideo_payload_endOfPack = 1'b0;
    if(when_Utils_l503_1) begin
      tmp_inputVideo_payload_endOfPack = 1'b1;
    end
  end

  always @(*) begin
    tmp_inputVideo_payload_endOfPack_1 = (tmp_inputVideo_payload_endOfPack_2 + tmp_tmp_inputVideo_payload_endOfPack_1);
    if(1'b0) begin
      tmp_inputVideo_payload_endOfPack_1 = 8'h0;
    end
  end

  assign tmp_when_Utils_l503 = (tmp_when_Utils_l503_4 == width);
  assign tmp_when_Utils_l503_1 = (tmp_when_Utils_l503_7 == height);
  assign inputVideo_valid = inputChannelSpilt_translated_m2sPipe_valid;
  assign inputChannelSpilt_translated_m2sPipe_ready = inputVideo_ready;
  assign inputVideo_payload_frame_line_pixel_0 = inputChannelSpilt_translated_m2sPipe_payload_0;
  assign inputVideo_payload_frame_line_pixel_1 = inputChannelSpilt_translated_m2sPipe_payload_1;
  assign inputVideo_payload_frame_line_pixel_2 = inputChannelSpilt_translated_m2sPipe_payload_2;
  assign inputVideo_payload_frame_line_pixel_3 = inputChannelSpilt_translated_m2sPipe_payload_3;
  assign inputVideo_payload_frame_line_pixel_4 = inputChannelSpilt_translated_m2sPipe_payload_4;
  assign inputVideo_payload_frame_line_pixel_5 = inputChannelSpilt_translated_m2sPipe_payload_5;
  assign inputVideo_payload_frame_line_pixel_6 = inputChannelSpilt_translated_m2sPipe_payload_6;
  assign inputVideo_payload_frame_line_pixel_7 = inputChannelSpilt_translated_m2sPipe_payload_7;
  assign inputVideo_payload_frame_line_pixel_8 = inputChannelSpilt_translated_m2sPipe_payload_8;
  assign inputVideo_payload_frame_line_pixel_9 = inputChannelSpilt_translated_m2sPipe_payload_9;
  assign inputVideo_payload_frame_line_pixel_10 = inputChannelSpilt_translated_m2sPipe_payload_10;
  assign inputVideo_payload_frame_line_pixel_11 = inputChannelSpilt_translated_m2sPipe_payload_11;
  assign inputVideo_payload_frame_line_pixel_12 = inputChannelSpilt_translated_m2sPipe_payload_12;
  assign inputVideo_payload_frame_line_pixel_13 = inputChannelSpilt_translated_m2sPipe_payload_13;
  assign inputVideo_payload_frame_line_pixel_14 = inputChannelSpilt_translated_m2sPipe_payload_14;
  assign inputVideo_payload_frame_line_pixel_15 = inputChannelSpilt_translated_m2sPipe_payload_15;
  assign inputVideo_payload_frame_line_endOfLine = tmp_when_Utils_l503;
  assign inputVideo_payload_frame_endOfFrame = tmp_when_Utils_l503_1;
  assign inputVideo_payload_endOfPack = (tmp_inputVideo_payload_endOfPack_2 == numberOfInputFrames);
  always @(*) begin
    tmp_io_select = 1'b0;
    if(weightsAdapted_fire) begin
      tmp_io_select = 1'b1;
    end
  end

  always @(*) begin
    tmp_io_select_1 = (tmp_io_select_2 + tmp_tmp_io_select_1);
    if(1'b0) begin
      tmp_io_select_1 = 3'b000;
    end
  end

  assign weightsAdapted_fire = (weightsAdapted_valid && weightsAdapted_ready);
  assign weightsAdapted_ready = streamDemux_2_io_input_ready;
  assign weights_fire = (weights_valid && weights_ready);
  always @(*) begin
    tmp_weights_ready = 1'b0;
    if(weights_fire) begin
      tmp_weights_ready = 1'b1;
    end
  end

  assign tmp_weights_ready_3 = (tmp_weights_ready_2 == 5'h11);
  assign tmp_1 = (tmp_weights_ready_3 && tmp_weights_ready);
  always @(*) begin
    if(tmp_1) begin
      tmp_weights_ready_1 = 5'h0;
    end else begin
      tmp_weights_ready_1 = (tmp_weights_ready_2 + tmp_tmp_weights_ready_1);
    end
    if(1'b0) begin
      tmp_weights_ready_1 = 5'h0;
    end
  end

  assign weights_fire_1 = (weights_valid && weights_ready);
  assign weightsAdapted_valid = (weights_valid && tmp_weights_ready_3);
  assign tmp_weightsAdapted_payload_0_0_0_0_1 = {weights_payload,tmp_weightsAdapted_payload_0_0_0_0};
  assign tmp_weightsAdapted_payload_0_0_0_0_2 = tmp_weightsAdapted_payload_0_0_0_0_1[1151 : 0];
  assign tmp_weightsAdapted_payload_0_0_0_0_3 = tmp_weightsAdapted_payload_0_0_0_0_2[383 : 0];
  assign tmp_weightsAdapted_payload_0_0_0_0_4 = tmp_weightsAdapted_payload_0_0_0_0_3[127 : 0];
  assign weightsAdapted_payload_0_0_0_0 = tmp_weightsAdapted_payload_0_0_0_0_4[7 : 0];
  assign weightsAdapted_payload_0_0_0_1 = tmp_weightsAdapted_payload_0_0_0_0_4[15 : 8];
  assign weightsAdapted_payload_0_0_0_2 = tmp_weightsAdapted_payload_0_0_0_0_4[23 : 16];
  assign weightsAdapted_payload_0_0_0_3 = tmp_weightsAdapted_payload_0_0_0_0_4[31 : 24];
  assign weightsAdapted_payload_0_0_0_4 = tmp_weightsAdapted_payload_0_0_0_0_4[39 : 32];
  assign weightsAdapted_payload_0_0_0_5 = tmp_weightsAdapted_payload_0_0_0_0_4[47 : 40];
  assign weightsAdapted_payload_0_0_0_6 = tmp_weightsAdapted_payload_0_0_0_0_4[55 : 48];
  assign weightsAdapted_payload_0_0_0_7 = tmp_weightsAdapted_payload_0_0_0_0_4[63 : 56];
  assign weightsAdapted_payload_0_0_0_8 = tmp_weightsAdapted_payload_0_0_0_0_4[71 : 64];
  assign weightsAdapted_payload_0_0_0_9 = tmp_weightsAdapted_payload_0_0_0_0_4[79 : 72];
  assign weightsAdapted_payload_0_0_0_10 = tmp_weightsAdapted_payload_0_0_0_0_4[87 : 80];
  assign weightsAdapted_payload_0_0_0_11 = tmp_weightsAdapted_payload_0_0_0_0_4[95 : 88];
  assign weightsAdapted_payload_0_0_0_12 = tmp_weightsAdapted_payload_0_0_0_0_4[103 : 96];
  assign weightsAdapted_payload_0_0_0_13 = tmp_weightsAdapted_payload_0_0_0_0_4[111 : 104];
  assign weightsAdapted_payload_0_0_0_14 = tmp_weightsAdapted_payload_0_0_0_0_4[119 : 112];
  assign weightsAdapted_payload_0_0_0_15 = tmp_weightsAdapted_payload_0_0_0_0_4[127 : 120];
  assign tmp_weightsAdapted_payload_0_0_1_0 = tmp_weightsAdapted_payload_0_0_0_0_3[255 : 128];
  assign weightsAdapted_payload_0_0_1_0 = tmp_weightsAdapted_payload_0_0_1_0[7 : 0];
  assign weightsAdapted_payload_0_0_1_1 = tmp_weightsAdapted_payload_0_0_1_0[15 : 8];
  assign weightsAdapted_payload_0_0_1_2 = tmp_weightsAdapted_payload_0_0_1_0[23 : 16];
  assign weightsAdapted_payload_0_0_1_3 = tmp_weightsAdapted_payload_0_0_1_0[31 : 24];
  assign weightsAdapted_payload_0_0_1_4 = tmp_weightsAdapted_payload_0_0_1_0[39 : 32];
  assign weightsAdapted_payload_0_0_1_5 = tmp_weightsAdapted_payload_0_0_1_0[47 : 40];
  assign weightsAdapted_payload_0_0_1_6 = tmp_weightsAdapted_payload_0_0_1_0[55 : 48];
  assign weightsAdapted_payload_0_0_1_7 = tmp_weightsAdapted_payload_0_0_1_0[63 : 56];
  assign weightsAdapted_payload_0_0_1_8 = tmp_weightsAdapted_payload_0_0_1_0[71 : 64];
  assign weightsAdapted_payload_0_0_1_9 = tmp_weightsAdapted_payload_0_0_1_0[79 : 72];
  assign weightsAdapted_payload_0_0_1_10 = tmp_weightsAdapted_payload_0_0_1_0[87 : 80];
  assign weightsAdapted_payload_0_0_1_11 = tmp_weightsAdapted_payload_0_0_1_0[95 : 88];
  assign weightsAdapted_payload_0_0_1_12 = tmp_weightsAdapted_payload_0_0_1_0[103 : 96];
  assign weightsAdapted_payload_0_0_1_13 = tmp_weightsAdapted_payload_0_0_1_0[111 : 104];
  assign weightsAdapted_payload_0_0_1_14 = tmp_weightsAdapted_payload_0_0_1_0[119 : 112];
  assign weightsAdapted_payload_0_0_1_15 = tmp_weightsAdapted_payload_0_0_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_0_0_2_0 = tmp_weightsAdapted_payload_0_0_0_0_3[383 : 256];
  assign weightsAdapted_payload_0_0_2_0 = tmp_weightsAdapted_payload_0_0_2_0[7 : 0];
  assign weightsAdapted_payload_0_0_2_1 = tmp_weightsAdapted_payload_0_0_2_0[15 : 8];
  assign weightsAdapted_payload_0_0_2_2 = tmp_weightsAdapted_payload_0_0_2_0[23 : 16];
  assign weightsAdapted_payload_0_0_2_3 = tmp_weightsAdapted_payload_0_0_2_0[31 : 24];
  assign weightsAdapted_payload_0_0_2_4 = tmp_weightsAdapted_payload_0_0_2_0[39 : 32];
  assign weightsAdapted_payload_0_0_2_5 = tmp_weightsAdapted_payload_0_0_2_0[47 : 40];
  assign weightsAdapted_payload_0_0_2_6 = tmp_weightsAdapted_payload_0_0_2_0[55 : 48];
  assign weightsAdapted_payload_0_0_2_7 = tmp_weightsAdapted_payload_0_0_2_0[63 : 56];
  assign weightsAdapted_payload_0_0_2_8 = tmp_weightsAdapted_payload_0_0_2_0[71 : 64];
  assign weightsAdapted_payload_0_0_2_9 = tmp_weightsAdapted_payload_0_0_2_0[79 : 72];
  assign weightsAdapted_payload_0_0_2_10 = tmp_weightsAdapted_payload_0_0_2_0[87 : 80];
  assign weightsAdapted_payload_0_0_2_11 = tmp_weightsAdapted_payload_0_0_2_0[95 : 88];
  assign weightsAdapted_payload_0_0_2_12 = tmp_weightsAdapted_payload_0_0_2_0[103 : 96];
  assign weightsAdapted_payload_0_0_2_13 = tmp_weightsAdapted_payload_0_0_2_0[111 : 104];
  assign weightsAdapted_payload_0_0_2_14 = tmp_weightsAdapted_payload_0_0_2_0[119 : 112];
  assign weightsAdapted_payload_0_0_2_15 = tmp_weightsAdapted_payload_0_0_2_0[127 : 120];
  assign tmp_weightsAdapted_payload_0_1_0_0 = tmp_weightsAdapted_payload_0_0_0_0_2[767 : 384];
  assign tmp_weightsAdapted_payload_0_1_0_0_1 = tmp_weightsAdapted_payload_0_1_0_0[127 : 0];
  assign weightsAdapted_payload_0_1_0_0 = tmp_weightsAdapted_payload_0_1_0_0_1[7 : 0];
  assign weightsAdapted_payload_0_1_0_1 = tmp_weightsAdapted_payload_0_1_0_0_1[15 : 8];
  assign weightsAdapted_payload_0_1_0_2 = tmp_weightsAdapted_payload_0_1_0_0_1[23 : 16];
  assign weightsAdapted_payload_0_1_0_3 = tmp_weightsAdapted_payload_0_1_0_0_1[31 : 24];
  assign weightsAdapted_payload_0_1_0_4 = tmp_weightsAdapted_payload_0_1_0_0_1[39 : 32];
  assign weightsAdapted_payload_0_1_0_5 = tmp_weightsAdapted_payload_0_1_0_0_1[47 : 40];
  assign weightsAdapted_payload_0_1_0_6 = tmp_weightsAdapted_payload_0_1_0_0_1[55 : 48];
  assign weightsAdapted_payload_0_1_0_7 = tmp_weightsAdapted_payload_0_1_0_0_1[63 : 56];
  assign weightsAdapted_payload_0_1_0_8 = tmp_weightsAdapted_payload_0_1_0_0_1[71 : 64];
  assign weightsAdapted_payload_0_1_0_9 = tmp_weightsAdapted_payload_0_1_0_0_1[79 : 72];
  assign weightsAdapted_payload_0_1_0_10 = tmp_weightsAdapted_payload_0_1_0_0_1[87 : 80];
  assign weightsAdapted_payload_0_1_0_11 = tmp_weightsAdapted_payload_0_1_0_0_1[95 : 88];
  assign weightsAdapted_payload_0_1_0_12 = tmp_weightsAdapted_payload_0_1_0_0_1[103 : 96];
  assign weightsAdapted_payload_0_1_0_13 = tmp_weightsAdapted_payload_0_1_0_0_1[111 : 104];
  assign weightsAdapted_payload_0_1_0_14 = tmp_weightsAdapted_payload_0_1_0_0_1[119 : 112];
  assign weightsAdapted_payload_0_1_0_15 = tmp_weightsAdapted_payload_0_1_0_0_1[127 : 120];
  assign tmp_weightsAdapted_payload_0_1_1_0 = tmp_weightsAdapted_payload_0_1_0_0[255 : 128];
  assign weightsAdapted_payload_0_1_1_0 = tmp_weightsAdapted_payload_0_1_1_0[7 : 0];
  assign weightsAdapted_payload_0_1_1_1 = tmp_weightsAdapted_payload_0_1_1_0[15 : 8];
  assign weightsAdapted_payload_0_1_1_2 = tmp_weightsAdapted_payload_0_1_1_0[23 : 16];
  assign weightsAdapted_payload_0_1_1_3 = tmp_weightsAdapted_payload_0_1_1_0[31 : 24];
  assign weightsAdapted_payload_0_1_1_4 = tmp_weightsAdapted_payload_0_1_1_0[39 : 32];
  assign weightsAdapted_payload_0_1_1_5 = tmp_weightsAdapted_payload_0_1_1_0[47 : 40];
  assign weightsAdapted_payload_0_1_1_6 = tmp_weightsAdapted_payload_0_1_1_0[55 : 48];
  assign weightsAdapted_payload_0_1_1_7 = tmp_weightsAdapted_payload_0_1_1_0[63 : 56];
  assign weightsAdapted_payload_0_1_1_8 = tmp_weightsAdapted_payload_0_1_1_0[71 : 64];
  assign weightsAdapted_payload_0_1_1_9 = tmp_weightsAdapted_payload_0_1_1_0[79 : 72];
  assign weightsAdapted_payload_0_1_1_10 = tmp_weightsAdapted_payload_0_1_1_0[87 : 80];
  assign weightsAdapted_payload_0_1_1_11 = tmp_weightsAdapted_payload_0_1_1_0[95 : 88];
  assign weightsAdapted_payload_0_1_1_12 = tmp_weightsAdapted_payload_0_1_1_0[103 : 96];
  assign weightsAdapted_payload_0_1_1_13 = tmp_weightsAdapted_payload_0_1_1_0[111 : 104];
  assign weightsAdapted_payload_0_1_1_14 = tmp_weightsAdapted_payload_0_1_1_0[119 : 112];
  assign weightsAdapted_payload_0_1_1_15 = tmp_weightsAdapted_payload_0_1_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_0_1_2_0 = tmp_weightsAdapted_payload_0_1_0_0[383 : 256];
  assign weightsAdapted_payload_0_1_2_0 = tmp_weightsAdapted_payload_0_1_2_0[7 : 0];
  assign weightsAdapted_payload_0_1_2_1 = tmp_weightsAdapted_payload_0_1_2_0[15 : 8];
  assign weightsAdapted_payload_0_1_2_2 = tmp_weightsAdapted_payload_0_1_2_0[23 : 16];
  assign weightsAdapted_payload_0_1_2_3 = tmp_weightsAdapted_payload_0_1_2_0[31 : 24];
  assign weightsAdapted_payload_0_1_2_4 = tmp_weightsAdapted_payload_0_1_2_0[39 : 32];
  assign weightsAdapted_payload_0_1_2_5 = tmp_weightsAdapted_payload_0_1_2_0[47 : 40];
  assign weightsAdapted_payload_0_1_2_6 = tmp_weightsAdapted_payload_0_1_2_0[55 : 48];
  assign weightsAdapted_payload_0_1_2_7 = tmp_weightsAdapted_payload_0_1_2_0[63 : 56];
  assign weightsAdapted_payload_0_1_2_8 = tmp_weightsAdapted_payload_0_1_2_0[71 : 64];
  assign weightsAdapted_payload_0_1_2_9 = tmp_weightsAdapted_payload_0_1_2_0[79 : 72];
  assign weightsAdapted_payload_0_1_2_10 = tmp_weightsAdapted_payload_0_1_2_0[87 : 80];
  assign weightsAdapted_payload_0_1_2_11 = tmp_weightsAdapted_payload_0_1_2_0[95 : 88];
  assign weightsAdapted_payload_0_1_2_12 = tmp_weightsAdapted_payload_0_1_2_0[103 : 96];
  assign weightsAdapted_payload_0_1_2_13 = tmp_weightsAdapted_payload_0_1_2_0[111 : 104];
  assign weightsAdapted_payload_0_1_2_14 = tmp_weightsAdapted_payload_0_1_2_0[119 : 112];
  assign weightsAdapted_payload_0_1_2_15 = tmp_weightsAdapted_payload_0_1_2_0[127 : 120];
  assign tmp_weightsAdapted_payload_0_2_0_0 = tmp_weightsAdapted_payload_0_0_0_0_2[1151 : 768];
  assign tmp_weightsAdapted_payload_0_2_0_0_1 = tmp_weightsAdapted_payload_0_2_0_0[127 : 0];
  assign weightsAdapted_payload_0_2_0_0 = tmp_weightsAdapted_payload_0_2_0_0_1[7 : 0];
  assign weightsAdapted_payload_0_2_0_1 = tmp_weightsAdapted_payload_0_2_0_0_1[15 : 8];
  assign weightsAdapted_payload_0_2_0_2 = tmp_weightsAdapted_payload_0_2_0_0_1[23 : 16];
  assign weightsAdapted_payload_0_2_0_3 = tmp_weightsAdapted_payload_0_2_0_0_1[31 : 24];
  assign weightsAdapted_payload_0_2_0_4 = tmp_weightsAdapted_payload_0_2_0_0_1[39 : 32];
  assign weightsAdapted_payload_0_2_0_5 = tmp_weightsAdapted_payload_0_2_0_0_1[47 : 40];
  assign weightsAdapted_payload_0_2_0_6 = tmp_weightsAdapted_payload_0_2_0_0_1[55 : 48];
  assign weightsAdapted_payload_0_2_0_7 = tmp_weightsAdapted_payload_0_2_0_0_1[63 : 56];
  assign weightsAdapted_payload_0_2_0_8 = tmp_weightsAdapted_payload_0_2_0_0_1[71 : 64];
  assign weightsAdapted_payload_0_2_0_9 = tmp_weightsAdapted_payload_0_2_0_0_1[79 : 72];
  assign weightsAdapted_payload_0_2_0_10 = tmp_weightsAdapted_payload_0_2_0_0_1[87 : 80];
  assign weightsAdapted_payload_0_2_0_11 = tmp_weightsAdapted_payload_0_2_0_0_1[95 : 88];
  assign weightsAdapted_payload_0_2_0_12 = tmp_weightsAdapted_payload_0_2_0_0_1[103 : 96];
  assign weightsAdapted_payload_0_2_0_13 = tmp_weightsAdapted_payload_0_2_0_0_1[111 : 104];
  assign weightsAdapted_payload_0_2_0_14 = tmp_weightsAdapted_payload_0_2_0_0_1[119 : 112];
  assign weightsAdapted_payload_0_2_0_15 = tmp_weightsAdapted_payload_0_2_0_0_1[127 : 120];
  assign tmp_weightsAdapted_payload_0_2_1_0 = tmp_weightsAdapted_payload_0_2_0_0[255 : 128];
  assign weightsAdapted_payload_0_2_1_0 = tmp_weightsAdapted_payload_0_2_1_0[7 : 0];
  assign weightsAdapted_payload_0_2_1_1 = tmp_weightsAdapted_payload_0_2_1_0[15 : 8];
  assign weightsAdapted_payload_0_2_1_2 = tmp_weightsAdapted_payload_0_2_1_0[23 : 16];
  assign weightsAdapted_payload_0_2_1_3 = tmp_weightsAdapted_payload_0_2_1_0[31 : 24];
  assign weightsAdapted_payload_0_2_1_4 = tmp_weightsAdapted_payload_0_2_1_0[39 : 32];
  assign weightsAdapted_payload_0_2_1_5 = tmp_weightsAdapted_payload_0_2_1_0[47 : 40];
  assign weightsAdapted_payload_0_2_1_6 = tmp_weightsAdapted_payload_0_2_1_0[55 : 48];
  assign weightsAdapted_payload_0_2_1_7 = tmp_weightsAdapted_payload_0_2_1_0[63 : 56];
  assign weightsAdapted_payload_0_2_1_8 = tmp_weightsAdapted_payload_0_2_1_0[71 : 64];
  assign weightsAdapted_payload_0_2_1_9 = tmp_weightsAdapted_payload_0_2_1_0[79 : 72];
  assign weightsAdapted_payload_0_2_1_10 = tmp_weightsAdapted_payload_0_2_1_0[87 : 80];
  assign weightsAdapted_payload_0_2_1_11 = tmp_weightsAdapted_payload_0_2_1_0[95 : 88];
  assign weightsAdapted_payload_0_2_1_12 = tmp_weightsAdapted_payload_0_2_1_0[103 : 96];
  assign weightsAdapted_payload_0_2_1_13 = tmp_weightsAdapted_payload_0_2_1_0[111 : 104];
  assign weightsAdapted_payload_0_2_1_14 = tmp_weightsAdapted_payload_0_2_1_0[119 : 112];
  assign weightsAdapted_payload_0_2_1_15 = tmp_weightsAdapted_payload_0_2_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_0_2_2_0 = tmp_weightsAdapted_payload_0_2_0_0[383 : 256];
  assign weightsAdapted_payload_0_2_2_0 = tmp_weightsAdapted_payload_0_2_2_0[7 : 0];
  assign weightsAdapted_payload_0_2_2_1 = tmp_weightsAdapted_payload_0_2_2_0[15 : 8];
  assign weightsAdapted_payload_0_2_2_2 = tmp_weightsAdapted_payload_0_2_2_0[23 : 16];
  assign weightsAdapted_payload_0_2_2_3 = tmp_weightsAdapted_payload_0_2_2_0[31 : 24];
  assign weightsAdapted_payload_0_2_2_4 = tmp_weightsAdapted_payload_0_2_2_0[39 : 32];
  assign weightsAdapted_payload_0_2_2_5 = tmp_weightsAdapted_payload_0_2_2_0[47 : 40];
  assign weightsAdapted_payload_0_2_2_6 = tmp_weightsAdapted_payload_0_2_2_0[55 : 48];
  assign weightsAdapted_payload_0_2_2_7 = tmp_weightsAdapted_payload_0_2_2_0[63 : 56];
  assign weightsAdapted_payload_0_2_2_8 = tmp_weightsAdapted_payload_0_2_2_0[71 : 64];
  assign weightsAdapted_payload_0_2_2_9 = tmp_weightsAdapted_payload_0_2_2_0[79 : 72];
  assign weightsAdapted_payload_0_2_2_10 = tmp_weightsAdapted_payload_0_2_2_0[87 : 80];
  assign weightsAdapted_payload_0_2_2_11 = tmp_weightsAdapted_payload_0_2_2_0[95 : 88];
  assign weightsAdapted_payload_0_2_2_12 = tmp_weightsAdapted_payload_0_2_2_0[103 : 96];
  assign weightsAdapted_payload_0_2_2_13 = tmp_weightsAdapted_payload_0_2_2_0[111 : 104];
  assign weightsAdapted_payload_0_2_2_14 = tmp_weightsAdapted_payload_0_2_2_0[119 : 112];
  assign weightsAdapted_payload_0_2_2_15 = tmp_weightsAdapted_payload_0_2_2_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_0_0_0 = tmp_weightsAdapted_payload_0_0_0_0_1[2303 : 1152];
  assign tmp_weightsAdapted_payload_1_0_0_0_1 = tmp_weightsAdapted_payload_1_0_0_0[383 : 0];
  assign tmp_weightsAdapted_payload_1_0_0_0_2 = tmp_weightsAdapted_payload_1_0_0_0_1[127 : 0];
  assign weightsAdapted_payload_1_0_0_0 = tmp_weightsAdapted_payload_1_0_0_0_2[7 : 0];
  assign weightsAdapted_payload_1_0_0_1 = tmp_weightsAdapted_payload_1_0_0_0_2[15 : 8];
  assign weightsAdapted_payload_1_0_0_2 = tmp_weightsAdapted_payload_1_0_0_0_2[23 : 16];
  assign weightsAdapted_payload_1_0_0_3 = tmp_weightsAdapted_payload_1_0_0_0_2[31 : 24];
  assign weightsAdapted_payload_1_0_0_4 = tmp_weightsAdapted_payload_1_0_0_0_2[39 : 32];
  assign weightsAdapted_payload_1_0_0_5 = tmp_weightsAdapted_payload_1_0_0_0_2[47 : 40];
  assign weightsAdapted_payload_1_0_0_6 = tmp_weightsAdapted_payload_1_0_0_0_2[55 : 48];
  assign weightsAdapted_payload_1_0_0_7 = tmp_weightsAdapted_payload_1_0_0_0_2[63 : 56];
  assign weightsAdapted_payload_1_0_0_8 = tmp_weightsAdapted_payload_1_0_0_0_2[71 : 64];
  assign weightsAdapted_payload_1_0_0_9 = tmp_weightsAdapted_payload_1_0_0_0_2[79 : 72];
  assign weightsAdapted_payload_1_0_0_10 = tmp_weightsAdapted_payload_1_0_0_0_2[87 : 80];
  assign weightsAdapted_payload_1_0_0_11 = tmp_weightsAdapted_payload_1_0_0_0_2[95 : 88];
  assign weightsAdapted_payload_1_0_0_12 = tmp_weightsAdapted_payload_1_0_0_0_2[103 : 96];
  assign weightsAdapted_payload_1_0_0_13 = tmp_weightsAdapted_payload_1_0_0_0_2[111 : 104];
  assign weightsAdapted_payload_1_0_0_14 = tmp_weightsAdapted_payload_1_0_0_0_2[119 : 112];
  assign weightsAdapted_payload_1_0_0_15 = tmp_weightsAdapted_payload_1_0_0_0_2[127 : 120];
  assign tmp_weightsAdapted_payload_1_0_1_0 = tmp_weightsAdapted_payload_1_0_0_0_1[255 : 128];
  assign weightsAdapted_payload_1_0_1_0 = tmp_weightsAdapted_payload_1_0_1_0[7 : 0];
  assign weightsAdapted_payload_1_0_1_1 = tmp_weightsAdapted_payload_1_0_1_0[15 : 8];
  assign weightsAdapted_payload_1_0_1_2 = tmp_weightsAdapted_payload_1_0_1_0[23 : 16];
  assign weightsAdapted_payload_1_0_1_3 = tmp_weightsAdapted_payload_1_0_1_0[31 : 24];
  assign weightsAdapted_payload_1_0_1_4 = tmp_weightsAdapted_payload_1_0_1_0[39 : 32];
  assign weightsAdapted_payload_1_0_1_5 = tmp_weightsAdapted_payload_1_0_1_0[47 : 40];
  assign weightsAdapted_payload_1_0_1_6 = tmp_weightsAdapted_payload_1_0_1_0[55 : 48];
  assign weightsAdapted_payload_1_0_1_7 = tmp_weightsAdapted_payload_1_0_1_0[63 : 56];
  assign weightsAdapted_payload_1_0_1_8 = tmp_weightsAdapted_payload_1_0_1_0[71 : 64];
  assign weightsAdapted_payload_1_0_1_9 = tmp_weightsAdapted_payload_1_0_1_0[79 : 72];
  assign weightsAdapted_payload_1_0_1_10 = tmp_weightsAdapted_payload_1_0_1_0[87 : 80];
  assign weightsAdapted_payload_1_0_1_11 = tmp_weightsAdapted_payload_1_0_1_0[95 : 88];
  assign weightsAdapted_payload_1_0_1_12 = tmp_weightsAdapted_payload_1_0_1_0[103 : 96];
  assign weightsAdapted_payload_1_0_1_13 = tmp_weightsAdapted_payload_1_0_1_0[111 : 104];
  assign weightsAdapted_payload_1_0_1_14 = tmp_weightsAdapted_payload_1_0_1_0[119 : 112];
  assign weightsAdapted_payload_1_0_1_15 = tmp_weightsAdapted_payload_1_0_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_0_2_0 = tmp_weightsAdapted_payload_1_0_0_0_1[383 : 256];
  assign weightsAdapted_payload_1_0_2_0 = tmp_weightsAdapted_payload_1_0_2_0[7 : 0];
  assign weightsAdapted_payload_1_0_2_1 = tmp_weightsAdapted_payload_1_0_2_0[15 : 8];
  assign weightsAdapted_payload_1_0_2_2 = tmp_weightsAdapted_payload_1_0_2_0[23 : 16];
  assign weightsAdapted_payload_1_0_2_3 = tmp_weightsAdapted_payload_1_0_2_0[31 : 24];
  assign weightsAdapted_payload_1_0_2_4 = tmp_weightsAdapted_payload_1_0_2_0[39 : 32];
  assign weightsAdapted_payload_1_0_2_5 = tmp_weightsAdapted_payload_1_0_2_0[47 : 40];
  assign weightsAdapted_payload_1_0_2_6 = tmp_weightsAdapted_payload_1_0_2_0[55 : 48];
  assign weightsAdapted_payload_1_0_2_7 = tmp_weightsAdapted_payload_1_0_2_0[63 : 56];
  assign weightsAdapted_payload_1_0_2_8 = tmp_weightsAdapted_payload_1_0_2_0[71 : 64];
  assign weightsAdapted_payload_1_0_2_9 = tmp_weightsAdapted_payload_1_0_2_0[79 : 72];
  assign weightsAdapted_payload_1_0_2_10 = tmp_weightsAdapted_payload_1_0_2_0[87 : 80];
  assign weightsAdapted_payload_1_0_2_11 = tmp_weightsAdapted_payload_1_0_2_0[95 : 88];
  assign weightsAdapted_payload_1_0_2_12 = tmp_weightsAdapted_payload_1_0_2_0[103 : 96];
  assign weightsAdapted_payload_1_0_2_13 = tmp_weightsAdapted_payload_1_0_2_0[111 : 104];
  assign weightsAdapted_payload_1_0_2_14 = tmp_weightsAdapted_payload_1_0_2_0[119 : 112];
  assign weightsAdapted_payload_1_0_2_15 = tmp_weightsAdapted_payload_1_0_2_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_1_0_0 = tmp_weightsAdapted_payload_1_0_0_0[767 : 384];
  assign tmp_weightsAdapted_payload_1_1_0_0_1 = tmp_weightsAdapted_payload_1_1_0_0[127 : 0];
  assign weightsAdapted_payload_1_1_0_0 = tmp_weightsAdapted_payload_1_1_0_0_1[7 : 0];
  assign weightsAdapted_payload_1_1_0_1 = tmp_weightsAdapted_payload_1_1_0_0_1[15 : 8];
  assign weightsAdapted_payload_1_1_0_2 = tmp_weightsAdapted_payload_1_1_0_0_1[23 : 16];
  assign weightsAdapted_payload_1_1_0_3 = tmp_weightsAdapted_payload_1_1_0_0_1[31 : 24];
  assign weightsAdapted_payload_1_1_0_4 = tmp_weightsAdapted_payload_1_1_0_0_1[39 : 32];
  assign weightsAdapted_payload_1_1_0_5 = tmp_weightsAdapted_payload_1_1_0_0_1[47 : 40];
  assign weightsAdapted_payload_1_1_0_6 = tmp_weightsAdapted_payload_1_1_0_0_1[55 : 48];
  assign weightsAdapted_payload_1_1_0_7 = tmp_weightsAdapted_payload_1_1_0_0_1[63 : 56];
  assign weightsAdapted_payload_1_1_0_8 = tmp_weightsAdapted_payload_1_1_0_0_1[71 : 64];
  assign weightsAdapted_payload_1_1_0_9 = tmp_weightsAdapted_payload_1_1_0_0_1[79 : 72];
  assign weightsAdapted_payload_1_1_0_10 = tmp_weightsAdapted_payload_1_1_0_0_1[87 : 80];
  assign weightsAdapted_payload_1_1_0_11 = tmp_weightsAdapted_payload_1_1_0_0_1[95 : 88];
  assign weightsAdapted_payload_1_1_0_12 = tmp_weightsAdapted_payload_1_1_0_0_1[103 : 96];
  assign weightsAdapted_payload_1_1_0_13 = tmp_weightsAdapted_payload_1_1_0_0_1[111 : 104];
  assign weightsAdapted_payload_1_1_0_14 = tmp_weightsAdapted_payload_1_1_0_0_1[119 : 112];
  assign weightsAdapted_payload_1_1_0_15 = tmp_weightsAdapted_payload_1_1_0_0_1[127 : 120];
  assign tmp_weightsAdapted_payload_1_1_1_0 = tmp_weightsAdapted_payload_1_1_0_0[255 : 128];
  assign weightsAdapted_payload_1_1_1_0 = tmp_weightsAdapted_payload_1_1_1_0[7 : 0];
  assign weightsAdapted_payload_1_1_1_1 = tmp_weightsAdapted_payload_1_1_1_0[15 : 8];
  assign weightsAdapted_payload_1_1_1_2 = tmp_weightsAdapted_payload_1_1_1_0[23 : 16];
  assign weightsAdapted_payload_1_1_1_3 = tmp_weightsAdapted_payload_1_1_1_0[31 : 24];
  assign weightsAdapted_payload_1_1_1_4 = tmp_weightsAdapted_payload_1_1_1_0[39 : 32];
  assign weightsAdapted_payload_1_1_1_5 = tmp_weightsAdapted_payload_1_1_1_0[47 : 40];
  assign weightsAdapted_payload_1_1_1_6 = tmp_weightsAdapted_payload_1_1_1_0[55 : 48];
  assign weightsAdapted_payload_1_1_1_7 = tmp_weightsAdapted_payload_1_1_1_0[63 : 56];
  assign weightsAdapted_payload_1_1_1_8 = tmp_weightsAdapted_payload_1_1_1_0[71 : 64];
  assign weightsAdapted_payload_1_1_1_9 = tmp_weightsAdapted_payload_1_1_1_0[79 : 72];
  assign weightsAdapted_payload_1_1_1_10 = tmp_weightsAdapted_payload_1_1_1_0[87 : 80];
  assign weightsAdapted_payload_1_1_1_11 = tmp_weightsAdapted_payload_1_1_1_0[95 : 88];
  assign weightsAdapted_payload_1_1_1_12 = tmp_weightsAdapted_payload_1_1_1_0[103 : 96];
  assign weightsAdapted_payload_1_1_1_13 = tmp_weightsAdapted_payload_1_1_1_0[111 : 104];
  assign weightsAdapted_payload_1_1_1_14 = tmp_weightsAdapted_payload_1_1_1_0[119 : 112];
  assign weightsAdapted_payload_1_1_1_15 = tmp_weightsAdapted_payload_1_1_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_1_2_0 = tmp_weightsAdapted_payload_1_1_0_0[383 : 256];
  assign weightsAdapted_payload_1_1_2_0 = tmp_weightsAdapted_payload_1_1_2_0[7 : 0];
  assign weightsAdapted_payload_1_1_2_1 = tmp_weightsAdapted_payload_1_1_2_0[15 : 8];
  assign weightsAdapted_payload_1_1_2_2 = tmp_weightsAdapted_payload_1_1_2_0[23 : 16];
  assign weightsAdapted_payload_1_1_2_3 = tmp_weightsAdapted_payload_1_1_2_0[31 : 24];
  assign weightsAdapted_payload_1_1_2_4 = tmp_weightsAdapted_payload_1_1_2_0[39 : 32];
  assign weightsAdapted_payload_1_1_2_5 = tmp_weightsAdapted_payload_1_1_2_0[47 : 40];
  assign weightsAdapted_payload_1_1_2_6 = tmp_weightsAdapted_payload_1_1_2_0[55 : 48];
  assign weightsAdapted_payload_1_1_2_7 = tmp_weightsAdapted_payload_1_1_2_0[63 : 56];
  assign weightsAdapted_payload_1_1_2_8 = tmp_weightsAdapted_payload_1_1_2_0[71 : 64];
  assign weightsAdapted_payload_1_1_2_9 = tmp_weightsAdapted_payload_1_1_2_0[79 : 72];
  assign weightsAdapted_payload_1_1_2_10 = tmp_weightsAdapted_payload_1_1_2_0[87 : 80];
  assign weightsAdapted_payload_1_1_2_11 = tmp_weightsAdapted_payload_1_1_2_0[95 : 88];
  assign weightsAdapted_payload_1_1_2_12 = tmp_weightsAdapted_payload_1_1_2_0[103 : 96];
  assign weightsAdapted_payload_1_1_2_13 = tmp_weightsAdapted_payload_1_1_2_0[111 : 104];
  assign weightsAdapted_payload_1_1_2_14 = tmp_weightsAdapted_payload_1_1_2_0[119 : 112];
  assign weightsAdapted_payload_1_1_2_15 = tmp_weightsAdapted_payload_1_1_2_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_2_0_0 = tmp_weightsAdapted_payload_1_0_0_0[1151 : 768];
  assign tmp_weightsAdapted_payload_1_2_0_0_1 = tmp_weightsAdapted_payload_1_2_0_0[127 : 0];
  assign weightsAdapted_payload_1_2_0_0 = tmp_weightsAdapted_payload_1_2_0_0_1[7 : 0];
  assign weightsAdapted_payload_1_2_0_1 = tmp_weightsAdapted_payload_1_2_0_0_1[15 : 8];
  assign weightsAdapted_payload_1_2_0_2 = tmp_weightsAdapted_payload_1_2_0_0_1[23 : 16];
  assign weightsAdapted_payload_1_2_0_3 = tmp_weightsAdapted_payload_1_2_0_0_1[31 : 24];
  assign weightsAdapted_payload_1_2_0_4 = tmp_weightsAdapted_payload_1_2_0_0_1[39 : 32];
  assign weightsAdapted_payload_1_2_0_5 = tmp_weightsAdapted_payload_1_2_0_0_1[47 : 40];
  assign weightsAdapted_payload_1_2_0_6 = tmp_weightsAdapted_payload_1_2_0_0_1[55 : 48];
  assign weightsAdapted_payload_1_2_0_7 = tmp_weightsAdapted_payload_1_2_0_0_1[63 : 56];
  assign weightsAdapted_payload_1_2_0_8 = tmp_weightsAdapted_payload_1_2_0_0_1[71 : 64];
  assign weightsAdapted_payload_1_2_0_9 = tmp_weightsAdapted_payload_1_2_0_0_1[79 : 72];
  assign weightsAdapted_payload_1_2_0_10 = tmp_weightsAdapted_payload_1_2_0_0_1[87 : 80];
  assign weightsAdapted_payload_1_2_0_11 = tmp_weightsAdapted_payload_1_2_0_0_1[95 : 88];
  assign weightsAdapted_payload_1_2_0_12 = tmp_weightsAdapted_payload_1_2_0_0_1[103 : 96];
  assign weightsAdapted_payload_1_2_0_13 = tmp_weightsAdapted_payload_1_2_0_0_1[111 : 104];
  assign weightsAdapted_payload_1_2_0_14 = tmp_weightsAdapted_payload_1_2_0_0_1[119 : 112];
  assign weightsAdapted_payload_1_2_0_15 = tmp_weightsAdapted_payload_1_2_0_0_1[127 : 120];
  assign tmp_weightsAdapted_payload_1_2_1_0 = tmp_weightsAdapted_payload_1_2_0_0[255 : 128];
  assign weightsAdapted_payload_1_2_1_0 = tmp_weightsAdapted_payload_1_2_1_0[7 : 0];
  assign weightsAdapted_payload_1_2_1_1 = tmp_weightsAdapted_payload_1_2_1_0[15 : 8];
  assign weightsAdapted_payload_1_2_1_2 = tmp_weightsAdapted_payload_1_2_1_0[23 : 16];
  assign weightsAdapted_payload_1_2_1_3 = tmp_weightsAdapted_payload_1_2_1_0[31 : 24];
  assign weightsAdapted_payload_1_2_1_4 = tmp_weightsAdapted_payload_1_2_1_0[39 : 32];
  assign weightsAdapted_payload_1_2_1_5 = tmp_weightsAdapted_payload_1_2_1_0[47 : 40];
  assign weightsAdapted_payload_1_2_1_6 = tmp_weightsAdapted_payload_1_2_1_0[55 : 48];
  assign weightsAdapted_payload_1_2_1_7 = tmp_weightsAdapted_payload_1_2_1_0[63 : 56];
  assign weightsAdapted_payload_1_2_1_8 = tmp_weightsAdapted_payload_1_2_1_0[71 : 64];
  assign weightsAdapted_payload_1_2_1_9 = tmp_weightsAdapted_payload_1_2_1_0[79 : 72];
  assign weightsAdapted_payload_1_2_1_10 = tmp_weightsAdapted_payload_1_2_1_0[87 : 80];
  assign weightsAdapted_payload_1_2_1_11 = tmp_weightsAdapted_payload_1_2_1_0[95 : 88];
  assign weightsAdapted_payload_1_2_1_12 = tmp_weightsAdapted_payload_1_2_1_0[103 : 96];
  assign weightsAdapted_payload_1_2_1_13 = tmp_weightsAdapted_payload_1_2_1_0[111 : 104];
  assign weightsAdapted_payload_1_2_1_14 = tmp_weightsAdapted_payload_1_2_1_0[119 : 112];
  assign weightsAdapted_payload_1_2_1_15 = tmp_weightsAdapted_payload_1_2_1_0[127 : 120];
  assign tmp_weightsAdapted_payload_1_2_2_0 = tmp_weightsAdapted_payload_1_2_0_0[383 : 256];
  assign weightsAdapted_payload_1_2_2_0 = tmp_weightsAdapted_payload_1_2_2_0[7 : 0];
  assign weightsAdapted_payload_1_2_2_1 = tmp_weightsAdapted_payload_1_2_2_0[15 : 8];
  assign weightsAdapted_payload_1_2_2_2 = tmp_weightsAdapted_payload_1_2_2_0[23 : 16];
  assign weightsAdapted_payload_1_2_2_3 = tmp_weightsAdapted_payload_1_2_2_0[31 : 24];
  assign weightsAdapted_payload_1_2_2_4 = tmp_weightsAdapted_payload_1_2_2_0[39 : 32];
  assign weightsAdapted_payload_1_2_2_5 = tmp_weightsAdapted_payload_1_2_2_0[47 : 40];
  assign weightsAdapted_payload_1_2_2_6 = tmp_weightsAdapted_payload_1_2_2_0[55 : 48];
  assign weightsAdapted_payload_1_2_2_7 = tmp_weightsAdapted_payload_1_2_2_0[63 : 56];
  assign weightsAdapted_payload_1_2_2_8 = tmp_weightsAdapted_payload_1_2_2_0[71 : 64];
  assign weightsAdapted_payload_1_2_2_9 = tmp_weightsAdapted_payload_1_2_2_0[79 : 72];
  assign weightsAdapted_payload_1_2_2_10 = tmp_weightsAdapted_payload_1_2_2_0[87 : 80];
  assign weightsAdapted_payload_1_2_2_11 = tmp_weightsAdapted_payload_1_2_2_0[95 : 88];
  assign weightsAdapted_payload_1_2_2_12 = tmp_weightsAdapted_payload_1_2_2_0[103 : 96];
  assign weightsAdapted_payload_1_2_2_13 = tmp_weightsAdapted_payload_1_2_2_0[111 : 104];
  assign weightsAdapted_payload_1_2_2_14 = tmp_weightsAdapted_payload_1_2_2_0[119 : 112];
  assign weightsAdapted_payload_1_2_2_15 = tmp_weightsAdapted_payload_1_2_2_0[127 : 120];
  assign weights_ready = (! ((! weightsAdapted_ready) && tmp_weights_ready_3));
  assign tmp_accOutputs_0_ready_1 = (tmp_accOutputs_0_ready && accOutputsJoin_ready);
  assign tmp_accOutputs_0_ready = (((((((accOutputs_0_valid && accOutputs_1_valid) && accOutputs_2_valid) && accOutputs_3_valid) && accOutputs_4_valid) && accOutputs_5_valid) && accOutputs_6_valid) && accOutputs_7_valid);
  assign accOutputs_0_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_1_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_2_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_3_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_4_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_5_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_6_ready = tmp_accOutputs_0_ready_1;
  assign accOutputs_7_ready = tmp_accOutputs_0_ready_1;
  assign accOutputsJoin_valid = tmp_accOutputs_0_ready;
  assign accOutputsJoin_payload_endOfPack = accOutputs_0_payload_endOfPack;
  assign accOutputsJoin_payload_frame_endOfFrame = accOutputs_0_payload_frame_endOfFrame;
  assign accOutputsJoin_payload_frame_line_endOfLine = accOutputs_0_payload_frame_line_endOfLine;
  assign tmp_accOutputsJoin_payload_frame_line_pixel_0 = {{accOutputs_7_payload_frame_line_pixel_1,accOutputs_7_payload_frame_line_pixel_0},{{accOutputs_6_payload_frame_line_pixel_1,accOutputs_6_payload_frame_line_pixel_0},{{accOutputs_5_payload_frame_line_pixel_1,accOutputs_5_payload_frame_line_pixel_0},{{accOutputs_4_payload_frame_line_pixel_1,accOutputs_4_payload_frame_line_pixel_0},{{accOutputs_3_payload_frame_line_pixel_1,accOutputs_3_payload_frame_line_pixel_0},{{accOutputs_2_payload_frame_line_pixel_1,accOutputs_2_payload_frame_line_pixel_0},{{accOutputs_1_payload_frame_line_pixel_1,accOutputs_1_payload_frame_line_pixel_0},{accOutputs_0_payload_frame_line_pixel_1,accOutputs_0_payload_frame_line_pixel_0}}}}}}}};
  assign accOutputsJoin_payload_frame_line_pixel_0 = tmp_accOutputsJoin_payload_frame_line_pixel_0[23 : 0];
  assign accOutputsJoin_payload_frame_line_pixel_1 = tmp_accOutputsJoin_payload_frame_line_pixel_0[47 : 24];
  assign accOutputsJoin_payload_frame_line_pixel_2 = tmp_accOutputsJoin_payload_frame_line_pixel_0[71 : 48];
  assign accOutputsJoin_payload_frame_line_pixel_3 = tmp_accOutputsJoin_payload_frame_line_pixel_0[95 : 72];
  assign accOutputsJoin_payload_frame_line_pixel_4 = tmp_accOutputsJoin_payload_frame_line_pixel_0[119 : 96];
  assign accOutputsJoin_payload_frame_line_pixel_5 = tmp_accOutputsJoin_payload_frame_line_pixel_0[143 : 120];
  assign accOutputsJoin_payload_frame_line_pixel_6 = tmp_accOutputsJoin_payload_frame_line_pixel_0[167 : 144];
  assign accOutputsJoin_payload_frame_line_pixel_7 = tmp_accOutputsJoin_payload_frame_line_pixel_0[191 : 168];
  assign accOutputsJoin_payload_frame_line_pixel_8 = tmp_accOutputsJoin_payload_frame_line_pixel_0[215 : 192];
  assign accOutputsJoin_payload_frame_line_pixel_9 = tmp_accOutputsJoin_payload_frame_line_pixel_0[239 : 216];
  assign accOutputsJoin_payload_frame_line_pixel_10 = tmp_accOutputsJoin_payload_frame_line_pixel_0[263 : 240];
  assign accOutputsJoin_payload_frame_line_pixel_11 = tmp_accOutputsJoin_payload_frame_line_pixel_0[287 : 264];
  assign accOutputsJoin_payload_frame_line_pixel_12 = tmp_accOutputsJoin_payload_frame_line_pixel_0[311 : 288];
  assign accOutputsJoin_payload_frame_line_pixel_13 = tmp_accOutputsJoin_payload_frame_line_pixel_0[335 : 312];
  assign accOutputsJoin_payload_frame_line_pixel_14 = tmp_accOutputsJoin_payload_frame_line_pixel_0[359 : 336];
  assign accOutputsJoin_payload_frame_line_pixel_15 = tmp_accOutputsJoin_payload_frame_line_pixel_0[383 : 360];
  assign accOutputsJoin_ready = eventM2sPipes_9_eventIn_ready;
  assign postProcessOutputs_payload_frame_line_pixel_0 = ($signed(scalerINT16_16_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_1 = ($signed(scalerINT16_17_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_2 = ($signed(scalerINT16_18_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_3 = ($signed(scalerINT16_19_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_4 = ($signed(scalerINT16_20_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_5 = ($signed(scalerINT16_21_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_6 = ($signed(scalerINT16_22_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_7 = ($signed(scalerINT16_23_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_8 = ($signed(scalerINT16_24_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_9 = ($signed(scalerINT16_25_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_10 = ($signed(scalerINT16_26_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_11 = ($signed(scalerINT16_27_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_12 = ($signed(scalerINT16_28_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_13 = ($signed(scalerINT16_29_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_14 = ($signed(scalerINT16_30_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_payload_frame_line_pixel_15 = ($signed(scalerINT16_31_dout) + $signed(outputZeroPoint));
  assign postProcessOutputs_valid = eventM2sPipes_9_eventOut_valid;
  assign postProcessOutputs_payload_endOfPack = tmp_postProcessOutputs_payload_endOfPack_5;
  assign postProcessOutputs_payload_frame_endOfFrame = tmp_postProcessOutputs_payload_frame_endOfFrame_5;
  assign postProcessOutputs_payload_frame_line_endOfLine = tmp_postProcessOutputs_payload_frame_line_endOfLine_5;
  assign postProcessOutputs_ready = streamDemux_3_io_input_ready;
  assign streamDemux_3_io_select = enablePooling;
  assign streamMux_1_io_select = enablePooling;
  assign streamMux_1_io_output_translated_valid = streamMux_1_io_output_valid;
  assign streamMux_1_io_output_translated_payload_0 = streamMux_1_io_output_payload_frame_line_pixel_0;
  assign streamMux_1_io_output_translated_payload_1 = streamMux_1_io_output_payload_frame_line_pixel_1;
  assign streamMux_1_io_output_translated_payload_2 = streamMux_1_io_output_payload_frame_line_pixel_2;
  assign streamMux_1_io_output_translated_payload_3 = streamMux_1_io_output_payload_frame_line_pixel_3;
  assign streamMux_1_io_output_translated_payload_4 = streamMux_1_io_output_payload_frame_line_pixel_4;
  assign streamMux_1_io_output_translated_payload_5 = streamMux_1_io_output_payload_frame_line_pixel_5;
  assign streamMux_1_io_output_translated_payload_6 = streamMux_1_io_output_payload_frame_line_pixel_6;
  assign streamMux_1_io_output_translated_payload_7 = streamMux_1_io_output_payload_frame_line_pixel_7;
  assign streamMux_1_io_output_translated_payload_8 = streamMux_1_io_output_payload_frame_line_pixel_8;
  assign streamMux_1_io_output_translated_payload_9 = streamMux_1_io_output_payload_frame_line_pixel_9;
  assign streamMux_1_io_output_translated_payload_10 = streamMux_1_io_output_payload_frame_line_pixel_10;
  assign streamMux_1_io_output_translated_payload_11 = streamMux_1_io_output_payload_frame_line_pixel_11;
  assign streamMux_1_io_output_translated_payload_12 = streamMux_1_io_output_payload_frame_line_pixel_12;
  assign streamMux_1_io_output_translated_payload_13 = streamMux_1_io_output_payload_frame_line_pixel_13;
  assign streamMux_1_io_output_translated_payload_14 = streamMux_1_io_output_payload_frame_line_pixel_14;
  assign streamMux_1_io_output_translated_payload_15 = streamMux_1_io_output_payload_frame_line_pixel_15;
  assign signalTrim_valid = streamMux_1_io_output_translated_valid;
  assign streamMux_1_io_output_translated_ready = signalTrim_ready;
  assign tmp_signalTrim_payload_0 = {streamMux_1_io_output_translated_payload_15,{streamMux_1_io_output_translated_payload_14,{streamMux_1_io_output_translated_payload_13,{streamMux_1_io_output_translated_payload_12,{streamMux_1_io_output_translated_payload_11,{streamMux_1_io_output_translated_payload_10,{streamMux_1_io_output_translated_payload_9,{streamMux_1_io_output_translated_payload_8,{streamMux_1_io_output_translated_payload_7,{streamMux_1_io_output_translated_payload_6,{streamMux_1_io_output_translated_payload_5,{streamMux_1_io_output_translated_payload_4,{streamMux_1_io_output_translated_payload_3,{streamMux_1_io_output_translated_payload_2,{streamMux_1_io_output_translated_payload_1,streamMux_1_io_output_translated_payload_0}}}}}}}}}}}}}}};
  assign signalTrim_payload_0 = tmp_signalTrim_payload_0[7 : 0];
  assign signalTrim_payload_1 = tmp_signalTrim_payload_0[15 : 8];
  assign signalTrim_payload_2 = tmp_signalTrim_payload_0[23 : 16];
  assign signalTrim_payload_3 = tmp_signalTrim_payload_0[31 : 24];
  assign signalTrim_payload_4 = tmp_signalTrim_payload_0[39 : 32];
  assign signalTrim_payload_5 = tmp_signalTrim_payload_0[47 : 40];
  assign signalTrim_payload_6 = tmp_signalTrim_payload_0[55 : 48];
  assign signalTrim_payload_7 = tmp_signalTrim_payload_0[63 : 56];
  assign signalTrim_payload_8 = tmp_signalTrim_payload_0[71 : 64];
  assign signalTrim_payload_9 = tmp_signalTrim_payload_0[79 : 72];
  assign signalTrim_payload_10 = tmp_signalTrim_payload_0[87 : 80];
  assign signalTrim_payload_11 = tmp_signalTrim_payload_0[95 : 88];
  assign signalTrim_payload_12 = tmp_signalTrim_payload_0[103 : 96];
  assign signalTrim_payload_13 = tmp_signalTrim_payload_0[111 : 104];
  assign signalTrim_payload_14 = tmp_signalTrim_payload_0[119 : 112];
  assign signalTrim_payload_15 = tmp_signalTrim_payload_0[127 : 120];
  assign tableAdapted_fire = (tableAdapted_valid && tableAdapted_ready);
  always @(*) begin
    tmp_funcTable_ready = 1'b0;
    if(tableAdapted_fire) begin
      tmp_funcTable_ready = 1'b1;
    end
  end

  assign tmp_funcTable_ready_3 = (tmp_funcTable_ready_2 == 4'b1111);
  always @(*) begin
    tmp_funcTable_ready_1 = (tmp_funcTable_ready_2 + tmp_tmp_funcTable_ready_1);
    if(1'b0) begin
      tmp_funcTable_ready_1 = 4'b0000;
    end
  end

  assign tableAdapted_valid = funcTable_valid;
  assign tmp_tableAdapted_payload = funcTable_payload;
  assign tableAdapted_payload = tmp_tableAdapted_payload_1;
  assign funcTable_ready = (tableAdapted_ready && tmp_funcTable_ready_3);
  assign tableAdapted_ready = table_1_newTable_ready;
  assign signalTrim_ready = table_1_index_ready;
  assign table_1_value_transmuted_valid = table_1_value_valid;
  assign table_1_value_transmuted_payload = {table_1_value_payload_15,{table_1_value_payload_14,{table_1_value_payload_13,{table_1_value_payload_12,{table_1_value_payload_11,{table_1_value_payload_10,{table_1_value_payload_9,{table_1_value_payload_8,{table_1_value_payload_7,{table_1_value_payload_6,{table_1_value_payload_5,{table_1_value_payload_4,{table_1_value_payload_3,{table_1_value_payload_2,{table_1_value_payload_1,table_1_value_payload_0}}}}}}}}}}}}}}};
  assign outputs_valid = table_1_value_transmuted_valid;
  assign table_1_value_transmuted_ready = outputs_ready;
  assign outputs_payload = table_1_value_transmuted_payload;
  assign inputVideo_ready = window_videoIn_ready;
  assign accOutputs_0_valid = unit_0_outputs_valid;
  assign accOutputs_0_payload_frame_line_pixel_0 = unit_0_outputs_payload_frame_line_pixel_0;
  assign accOutputs_0_payload_frame_line_pixel_1 = unit_0_outputs_payload_frame_line_pixel_1;
  assign accOutputs_0_payload_frame_line_endOfLine = unit_0_outputs_payload_frame_line_endOfLine;
  assign accOutputs_0_payload_frame_endOfFrame = unit_0_outputs_payload_frame_endOfFrame;
  assign accOutputs_0_payload_endOfPack = unit_0_outputs_payload_endOfPack;
  assign accOutputs_1_valid = unit_1_outputs_valid;
  assign accOutputs_1_payload_frame_line_pixel_0 = unit_1_outputs_payload_frame_line_pixel_0;
  assign accOutputs_1_payload_frame_line_pixel_1 = unit_1_outputs_payload_frame_line_pixel_1;
  assign accOutputs_1_payload_frame_line_endOfLine = unit_1_outputs_payload_frame_line_endOfLine;
  assign accOutputs_1_payload_frame_endOfFrame = unit_1_outputs_payload_frame_endOfFrame;
  assign accOutputs_1_payload_endOfPack = unit_1_outputs_payload_endOfPack;
  assign accOutputs_2_valid = unit_2_outputs_valid;
  assign accOutputs_2_payload_frame_line_pixel_0 = unit_2_outputs_payload_frame_line_pixel_0;
  assign accOutputs_2_payload_frame_line_pixel_1 = unit_2_outputs_payload_frame_line_pixel_1;
  assign accOutputs_2_payload_frame_line_endOfLine = unit_2_outputs_payload_frame_line_endOfLine;
  assign accOutputs_2_payload_frame_endOfFrame = unit_2_outputs_payload_frame_endOfFrame;
  assign accOutputs_2_payload_endOfPack = unit_2_outputs_payload_endOfPack;
  assign accOutputs_3_valid = unit_3_outputs_valid;
  assign accOutputs_3_payload_frame_line_pixel_0 = unit_3_outputs_payload_frame_line_pixel_0;
  assign accOutputs_3_payload_frame_line_pixel_1 = unit_3_outputs_payload_frame_line_pixel_1;
  assign accOutputs_3_payload_frame_line_endOfLine = unit_3_outputs_payload_frame_line_endOfLine;
  assign accOutputs_3_payload_frame_endOfFrame = unit_3_outputs_payload_frame_endOfFrame;
  assign accOutputs_3_payload_endOfPack = unit_3_outputs_payload_endOfPack;
  assign accOutputs_4_valid = unit_4_outputs_valid;
  assign accOutputs_4_payload_frame_line_pixel_0 = unit_4_outputs_payload_frame_line_pixel_0;
  assign accOutputs_4_payload_frame_line_pixel_1 = unit_4_outputs_payload_frame_line_pixel_1;
  assign accOutputs_4_payload_frame_line_endOfLine = unit_4_outputs_payload_frame_line_endOfLine;
  assign accOutputs_4_payload_frame_endOfFrame = unit_4_outputs_payload_frame_endOfFrame;
  assign accOutputs_4_payload_endOfPack = unit_4_outputs_payload_endOfPack;
  assign accOutputs_5_valid = unit_5_outputs_valid;
  assign accOutputs_5_payload_frame_line_pixel_0 = unit_5_outputs_payload_frame_line_pixel_0;
  assign accOutputs_5_payload_frame_line_pixel_1 = unit_5_outputs_payload_frame_line_pixel_1;
  assign accOutputs_5_payload_frame_line_endOfLine = unit_5_outputs_payload_frame_line_endOfLine;
  assign accOutputs_5_payload_frame_endOfFrame = unit_5_outputs_payload_frame_endOfFrame;
  assign accOutputs_5_payload_endOfPack = unit_5_outputs_payload_endOfPack;
  assign accOutputs_6_valid = unit_6_outputs_valid;
  assign accOutputs_6_payload_frame_line_pixel_0 = unit_6_outputs_payload_frame_line_pixel_0;
  assign accOutputs_6_payload_frame_line_pixel_1 = unit_6_outputs_payload_frame_line_pixel_1;
  assign accOutputs_6_payload_frame_line_endOfLine = unit_6_outputs_payload_frame_line_endOfLine;
  assign accOutputs_6_payload_frame_endOfFrame = unit_6_outputs_payload_frame_endOfFrame;
  assign accOutputs_6_payload_endOfPack = unit_6_outputs_payload_endOfPack;
  assign accOutputs_7_valid = unit_7_outputs_valid;
  assign accOutputs_7_payload_frame_line_pixel_0 = unit_7_outputs_payload_frame_line_pixel_0;
  assign accOutputs_7_payload_frame_line_pixel_1 = unit_7_outputs_payload_frame_line_pixel_1;
  assign accOutputs_7_payload_frame_line_endOfLine = unit_7_outputs_payload_frame_line_endOfLine;
  assign accOutputs_7_payload_frame_endOfFrame = unit_7_outputs_payload_frame_endOfFrame;
  assign accOutputs_7_payload_endOfPack = unit_7_outputs_payload_endOfPack;
  always @(posedge clk) begin
    if(reset) begin
      inputChannelSpilt_translated_rValid <= 1'b0;
      tmp_when_Utils_l503_4 <= 9'h0;
      tmp_when_Utils_l503_7 <= 9'h0;
      tmp_inputVideo_payload_endOfPack_2 <= 8'h0;
      tmp_io_select_2 <= 3'b000;
      tmp_weights_ready_2 <= 5'h0;
      tmp_funcTable_ready_2 <= 4'b0000;
    end else begin
      if(inputChannelSpilt_translated_ready) begin
        inputChannelSpilt_translated_rValid <= inputChannelSpilt_translated_valid;
      end
      tmp_when_Utils_l503_4 <= tmp_when_Utils_l503_3;
      tmp_when_Utils_l503_7 <= tmp_when_Utils_l503_6;
      tmp_inputVideo_payload_endOfPack_2 <= tmp_inputVideo_payload_endOfPack_1;
      tmp_io_select_2 <= tmp_io_select_1;
      tmp_weights_ready_2 <= tmp_weights_ready_1;
      tmp_funcTable_ready_2 <= tmp_funcTable_ready_1;
    end
  end

  always @(posedge clk) begin
    if(inputChannelSpilt_translated_ready) begin
      inputChannelSpilt_translated_rData_0 <= inputChannelSpilt_translated_payload_0;
      inputChannelSpilt_translated_rData_1 <= inputChannelSpilt_translated_payload_1;
      inputChannelSpilt_translated_rData_2 <= inputChannelSpilt_translated_payload_2;
      inputChannelSpilt_translated_rData_3 <= inputChannelSpilt_translated_payload_3;
      inputChannelSpilt_translated_rData_4 <= inputChannelSpilt_translated_payload_4;
      inputChannelSpilt_translated_rData_5 <= inputChannelSpilt_translated_payload_5;
      inputChannelSpilt_translated_rData_6 <= inputChannelSpilt_translated_payload_6;
      inputChannelSpilt_translated_rData_7 <= inputChannelSpilt_translated_payload_7;
      inputChannelSpilt_translated_rData_8 <= inputChannelSpilt_translated_payload_8;
      inputChannelSpilt_translated_rData_9 <= inputChannelSpilt_translated_payload_9;
      inputChannelSpilt_translated_rData_10 <= inputChannelSpilt_translated_payload_10;
      inputChannelSpilt_translated_rData_11 <= inputChannelSpilt_translated_payload_11;
      inputChannelSpilt_translated_rData_12 <= inputChannelSpilt_translated_payload_12;
      inputChannelSpilt_translated_rData_13 <= inputChannelSpilt_translated_payload_13;
      inputChannelSpilt_translated_rData_14 <= inputChannelSpilt_translated_payload_14;
      inputChannelSpilt_translated_rData_15 <= inputChannelSpilt_translated_payload_15;
    end
    if(weights_fire_1) begin
      tmp_weightsAdapted_payload_0_0_0_0 <= {weights_payload,tmp_tmp_weightsAdapted_payload_0_0_0_0};
    end
    if(eventM2sPipes_9_CEs_0) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine <= accOutputsJoin_payload_frame_line_endOfLine;
      tmp_postProcessOutputs_payload_frame_endOfFrame <= accOutputsJoin_payload_frame_endOfFrame;
      tmp_postProcessOutputs_payload_endOfPack <= accOutputsJoin_payload_endOfPack;
    end
    if(eventM2sPipes_9_CEs_1) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine_1 <= tmp_postProcessOutputs_payload_frame_line_endOfLine;
      tmp_postProcessOutputs_payload_frame_endOfFrame_1 <= tmp_postProcessOutputs_payload_frame_endOfFrame;
      tmp_postProcessOutputs_payload_endOfPack_1 <= tmp_postProcessOutputs_payload_endOfPack;
    end
    if(eventM2sPipes_9_CEs_2) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine_2 <= tmp_postProcessOutputs_payload_frame_line_endOfLine_1;
      tmp_postProcessOutputs_payload_frame_endOfFrame_2 <= tmp_postProcessOutputs_payload_frame_endOfFrame_1;
      tmp_postProcessOutputs_payload_endOfPack_2 <= tmp_postProcessOutputs_payload_endOfPack_1;
    end
    if(eventM2sPipes_9_CEs_3) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine_3 <= tmp_postProcessOutputs_payload_frame_line_endOfLine_2;
      tmp_postProcessOutputs_payload_frame_endOfFrame_3 <= tmp_postProcessOutputs_payload_frame_endOfFrame_2;
      tmp_postProcessOutputs_payload_endOfPack_3 <= tmp_postProcessOutputs_payload_endOfPack_2;
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine_4 <= tmp_postProcessOutputs_payload_frame_line_endOfLine_3;
      tmp_postProcessOutputs_payload_frame_endOfFrame_4 <= tmp_postProcessOutputs_payload_frame_endOfFrame_3;
      tmp_postProcessOutputs_payload_endOfPack_4 <= tmp_postProcessOutputs_payload_endOfPack_3;
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postProcessOutputs_payload_frame_line_endOfLine_5 <= tmp_postProcessOutputs_payload_frame_line_endOfLine_4;
      tmp_postProcessOutputs_payload_frame_endOfFrame_5 <= tmp_postProcessOutputs_payload_frame_endOfFrame_4;
      tmp_postProcessOutputs_payload_endOfPack_5 <= tmp_postProcessOutputs_payload_endOfPack_4;
    end
  end


endmodule

module StreamMux (
  input      [0:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_0,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_1,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_2,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_3,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_4,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_5,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_6,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_7,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_8,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_9,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_10,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_11,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_12,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_13,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_14,
  input      [7:0]    io_inputs_0_payload_frame_line_pixel_15,
  input               io_inputs_0_payload_frame_line_endOfLine,
  input               io_inputs_0_payload_frame_endOfFrame,
  input               io_inputs_0_payload_endOfPack,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_0,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_1,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_2,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_3,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_4,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_5,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_6,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_7,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_8,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_9,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_10,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_11,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_12,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_13,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_14,
  input      [7:0]    io_inputs_1_payload_frame_line_pixel_15,
  input               io_inputs_1_payload_frame_line_endOfLine,
  input               io_inputs_1_payload_frame_endOfFrame,
  input               io_inputs_1_payload_endOfPack,
  output              io_output_valid,
  input               io_output_ready,
  output     [7:0]    io_output_payload_frame_line_pixel_0,
  output     [7:0]    io_output_payload_frame_line_pixel_1,
  output     [7:0]    io_output_payload_frame_line_pixel_2,
  output     [7:0]    io_output_payload_frame_line_pixel_3,
  output     [7:0]    io_output_payload_frame_line_pixel_4,
  output     [7:0]    io_output_payload_frame_line_pixel_5,
  output     [7:0]    io_output_payload_frame_line_pixel_6,
  output     [7:0]    io_output_payload_frame_line_pixel_7,
  output     [7:0]    io_output_payload_frame_line_pixel_8,
  output     [7:0]    io_output_payload_frame_line_pixel_9,
  output     [7:0]    io_output_payload_frame_line_pixel_10,
  output     [7:0]    io_output_payload_frame_line_pixel_11,
  output     [7:0]    io_output_payload_frame_line_pixel_12,
  output     [7:0]    io_output_payload_frame_line_pixel_13,
  output     [7:0]    io_output_payload_frame_line_pixel_14,
  output     [7:0]    io_output_payload_frame_line_pixel_15,
  output              io_output_payload_frame_line_endOfLine,
  output              io_output_payload_frame_endOfFrame,
  output              io_output_payload_endOfPack
);

  reg                 tmp_io_output_valid;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_0;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_1;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_2;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_3;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_4;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_5;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_6;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_7;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_8;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_9;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_10;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_11;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_12;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_13;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_14;
  reg        [7:0]    tmp_io_output_payload_frame_line_pixel_15;
  reg                 tmp_io_output_payload_frame_line_endOfLine;
  reg                 tmp_io_output_payload_frame_endOfFrame;
  reg                 tmp_io_output_payload_endOfPack;

  always @(*) begin
    case(io_select)
      1'b0 : begin
        tmp_io_output_valid = io_inputs_0_valid;
        tmp_io_output_payload_frame_line_pixel_0 = io_inputs_0_payload_frame_line_pixel_0;
        tmp_io_output_payload_frame_line_pixel_1 = io_inputs_0_payload_frame_line_pixel_1;
        tmp_io_output_payload_frame_line_pixel_2 = io_inputs_0_payload_frame_line_pixel_2;
        tmp_io_output_payload_frame_line_pixel_3 = io_inputs_0_payload_frame_line_pixel_3;
        tmp_io_output_payload_frame_line_pixel_4 = io_inputs_0_payload_frame_line_pixel_4;
        tmp_io_output_payload_frame_line_pixel_5 = io_inputs_0_payload_frame_line_pixel_5;
        tmp_io_output_payload_frame_line_pixel_6 = io_inputs_0_payload_frame_line_pixel_6;
        tmp_io_output_payload_frame_line_pixel_7 = io_inputs_0_payload_frame_line_pixel_7;
        tmp_io_output_payload_frame_line_pixel_8 = io_inputs_0_payload_frame_line_pixel_8;
        tmp_io_output_payload_frame_line_pixel_9 = io_inputs_0_payload_frame_line_pixel_9;
        tmp_io_output_payload_frame_line_pixel_10 = io_inputs_0_payload_frame_line_pixel_10;
        tmp_io_output_payload_frame_line_pixel_11 = io_inputs_0_payload_frame_line_pixel_11;
        tmp_io_output_payload_frame_line_pixel_12 = io_inputs_0_payload_frame_line_pixel_12;
        tmp_io_output_payload_frame_line_pixel_13 = io_inputs_0_payload_frame_line_pixel_13;
        tmp_io_output_payload_frame_line_pixel_14 = io_inputs_0_payload_frame_line_pixel_14;
        tmp_io_output_payload_frame_line_pixel_15 = io_inputs_0_payload_frame_line_pixel_15;
        tmp_io_output_payload_frame_line_endOfLine = io_inputs_0_payload_frame_line_endOfLine;
        tmp_io_output_payload_frame_endOfFrame = io_inputs_0_payload_frame_endOfFrame;
        tmp_io_output_payload_endOfPack = io_inputs_0_payload_endOfPack;
      end
      default : begin
        tmp_io_output_valid = io_inputs_1_valid;
        tmp_io_output_payload_frame_line_pixel_0 = io_inputs_1_payload_frame_line_pixel_0;
        tmp_io_output_payload_frame_line_pixel_1 = io_inputs_1_payload_frame_line_pixel_1;
        tmp_io_output_payload_frame_line_pixel_2 = io_inputs_1_payload_frame_line_pixel_2;
        tmp_io_output_payload_frame_line_pixel_3 = io_inputs_1_payload_frame_line_pixel_3;
        tmp_io_output_payload_frame_line_pixel_4 = io_inputs_1_payload_frame_line_pixel_4;
        tmp_io_output_payload_frame_line_pixel_5 = io_inputs_1_payload_frame_line_pixel_5;
        tmp_io_output_payload_frame_line_pixel_6 = io_inputs_1_payload_frame_line_pixel_6;
        tmp_io_output_payload_frame_line_pixel_7 = io_inputs_1_payload_frame_line_pixel_7;
        tmp_io_output_payload_frame_line_pixel_8 = io_inputs_1_payload_frame_line_pixel_8;
        tmp_io_output_payload_frame_line_pixel_9 = io_inputs_1_payload_frame_line_pixel_9;
        tmp_io_output_payload_frame_line_pixel_10 = io_inputs_1_payload_frame_line_pixel_10;
        tmp_io_output_payload_frame_line_pixel_11 = io_inputs_1_payload_frame_line_pixel_11;
        tmp_io_output_payload_frame_line_pixel_12 = io_inputs_1_payload_frame_line_pixel_12;
        tmp_io_output_payload_frame_line_pixel_13 = io_inputs_1_payload_frame_line_pixel_13;
        tmp_io_output_payload_frame_line_pixel_14 = io_inputs_1_payload_frame_line_pixel_14;
        tmp_io_output_payload_frame_line_pixel_15 = io_inputs_1_payload_frame_line_pixel_15;
        tmp_io_output_payload_frame_line_endOfLine = io_inputs_1_payload_frame_line_endOfLine;
        tmp_io_output_payload_frame_endOfFrame = io_inputs_1_payload_frame_endOfFrame;
        tmp_io_output_payload_endOfPack = io_inputs_1_payload_endOfPack;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 1'b0) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 1'b1) && io_output_ready);
  assign io_output_valid = tmp_io_output_valid;
  assign io_output_payload_frame_line_pixel_0 = tmp_io_output_payload_frame_line_pixel_0;
  assign io_output_payload_frame_line_pixel_1 = tmp_io_output_payload_frame_line_pixel_1;
  assign io_output_payload_frame_line_pixel_2 = tmp_io_output_payload_frame_line_pixel_2;
  assign io_output_payload_frame_line_pixel_3 = tmp_io_output_payload_frame_line_pixel_3;
  assign io_output_payload_frame_line_pixel_4 = tmp_io_output_payload_frame_line_pixel_4;
  assign io_output_payload_frame_line_pixel_5 = tmp_io_output_payload_frame_line_pixel_5;
  assign io_output_payload_frame_line_pixel_6 = tmp_io_output_payload_frame_line_pixel_6;
  assign io_output_payload_frame_line_pixel_7 = tmp_io_output_payload_frame_line_pixel_7;
  assign io_output_payload_frame_line_pixel_8 = tmp_io_output_payload_frame_line_pixel_8;
  assign io_output_payload_frame_line_pixel_9 = tmp_io_output_payload_frame_line_pixel_9;
  assign io_output_payload_frame_line_pixel_10 = tmp_io_output_payload_frame_line_pixel_10;
  assign io_output_payload_frame_line_pixel_11 = tmp_io_output_payload_frame_line_pixel_11;
  assign io_output_payload_frame_line_pixel_12 = tmp_io_output_payload_frame_line_pixel_12;
  assign io_output_payload_frame_line_pixel_13 = tmp_io_output_payload_frame_line_pixel_13;
  assign io_output_payload_frame_line_pixel_14 = tmp_io_output_payload_frame_line_pixel_14;
  assign io_output_payload_frame_line_pixel_15 = tmp_io_output_payload_frame_line_pixel_15;
  assign io_output_payload_frame_line_endOfLine = tmp_io_output_payload_frame_line_endOfLine;
  assign io_output_payload_frame_endOfFrame = tmp_io_output_payload_frame_endOfFrame;
  assign io_output_payload_endOfPack = tmp_io_output_payload_endOfPack;

endmodule

module StreamDemux_1 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_frame_line_pixel_0,
  input      [7:0]    io_input_payload_frame_line_pixel_1,
  input      [7:0]    io_input_payload_frame_line_pixel_2,
  input      [7:0]    io_input_payload_frame_line_pixel_3,
  input      [7:0]    io_input_payload_frame_line_pixel_4,
  input      [7:0]    io_input_payload_frame_line_pixel_5,
  input      [7:0]    io_input_payload_frame_line_pixel_6,
  input      [7:0]    io_input_payload_frame_line_pixel_7,
  input      [7:0]    io_input_payload_frame_line_pixel_8,
  input      [7:0]    io_input_payload_frame_line_pixel_9,
  input      [7:0]    io_input_payload_frame_line_pixel_10,
  input      [7:0]    io_input_payload_frame_line_pixel_11,
  input      [7:0]    io_input_payload_frame_line_pixel_12,
  input      [7:0]    io_input_payload_frame_line_pixel_13,
  input      [7:0]    io_input_payload_frame_line_pixel_14,
  input      [7:0]    io_input_payload_frame_line_pixel_15,
  input               io_input_payload_frame_line_endOfLine,
  input               io_input_payload_frame_endOfFrame,
  input               io_input_payload_endOfPack,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_15,
  output              io_outputs_0_payload_frame_line_endOfLine,
  output              io_outputs_0_payload_frame_endOfFrame,
  output              io_outputs_0_payload_endOfPack,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_15,
  output              io_outputs_1_payload_frame_line_endOfLine,
  output              io_outputs_1_payload_frame_endOfFrame,
  output              io_outputs_1_payload_endOfPack
);

  wire                when_Stream_l764;
  wire                when_Stream_l764_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l764) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l764_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_frame_line_pixel_0 = io_input_payload_frame_line_pixel_0;
  assign io_outputs_0_payload_frame_line_pixel_1 = io_input_payload_frame_line_pixel_1;
  assign io_outputs_0_payload_frame_line_pixel_2 = io_input_payload_frame_line_pixel_2;
  assign io_outputs_0_payload_frame_line_pixel_3 = io_input_payload_frame_line_pixel_3;
  assign io_outputs_0_payload_frame_line_pixel_4 = io_input_payload_frame_line_pixel_4;
  assign io_outputs_0_payload_frame_line_pixel_5 = io_input_payload_frame_line_pixel_5;
  assign io_outputs_0_payload_frame_line_pixel_6 = io_input_payload_frame_line_pixel_6;
  assign io_outputs_0_payload_frame_line_pixel_7 = io_input_payload_frame_line_pixel_7;
  assign io_outputs_0_payload_frame_line_pixel_8 = io_input_payload_frame_line_pixel_8;
  assign io_outputs_0_payload_frame_line_pixel_9 = io_input_payload_frame_line_pixel_9;
  assign io_outputs_0_payload_frame_line_pixel_10 = io_input_payload_frame_line_pixel_10;
  assign io_outputs_0_payload_frame_line_pixel_11 = io_input_payload_frame_line_pixel_11;
  assign io_outputs_0_payload_frame_line_pixel_12 = io_input_payload_frame_line_pixel_12;
  assign io_outputs_0_payload_frame_line_pixel_13 = io_input_payload_frame_line_pixel_13;
  assign io_outputs_0_payload_frame_line_pixel_14 = io_input_payload_frame_line_pixel_14;
  assign io_outputs_0_payload_frame_line_pixel_15 = io_input_payload_frame_line_pixel_15;
  assign io_outputs_0_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_0_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_0_payload_endOfPack = io_input_payload_endOfPack;
  assign when_Stream_l764 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l764) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_frame_line_pixel_0 = io_input_payload_frame_line_pixel_0;
  assign io_outputs_1_payload_frame_line_pixel_1 = io_input_payload_frame_line_pixel_1;
  assign io_outputs_1_payload_frame_line_pixel_2 = io_input_payload_frame_line_pixel_2;
  assign io_outputs_1_payload_frame_line_pixel_3 = io_input_payload_frame_line_pixel_3;
  assign io_outputs_1_payload_frame_line_pixel_4 = io_input_payload_frame_line_pixel_4;
  assign io_outputs_1_payload_frame_line_pixel_5 = io_input_payload_frame_line_pixel_5;
  assign io_outputs_1_payload_frame_line_pixel_6 = io_input_payload_frame_line_pixel_6;
  assign io_outputs_1_payload_frame_line_pixel_7 = io_input_payload_frame_line_pixel_7;
  assign io_outputs_1_payload_frame_line_pixel_8 = io_input_payload_frame_line_pixel_8;
  assign io_outputs_1_payload_frame_line_pixel_9 = io_input_payload_frame_line_pixel_9;
  assign io_outputs_1_payload_frame_line_pixel_10 = io_input_payload_frame_line_pixel_10;
  assign io_outputs_1_payload_frame_line_pixel_11 = io_input_payload_frame_line_pixel_11;
  assign io_outputs_1_payload_frame_line_pixel_12 = io_input_payload_frame_line_pixel_12;
  assign io_outputs_1_payload_frame_line_pixel_13 = io_input_payload_frame_line_pixel_13;
  assign io_outputs_1_payload_frame_line_pixel_14 = io_input_payload_frame_line_pixel_14;
  assign io_outputs_1_payload_frame_line_pixel_15 = io_input_payload_frame_line_pixel_15;
  assign io_outputs_1_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_1_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_1_payload_endOfPack = io_input_payload_endOfPack;
  assign when_Stream_l764_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l764_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

//ScalerINT16 replaced by ScalerINT16

module ScalerINT16 (
  input      [15:0]   scalerBase,
  input      [5:0]    scalerExpr,
  input               CEs_0,
  input               CEs_1,
  input               CEs_2,
  input               CEs_3,
  input               CEs_4,
  input               CEs_5,
  input      [23:0]   din,
  output     [7:0]    dout,
  input               clk,
  input               reset
);

  wire       [29:0]   mult_A;
  wire       [17:0]   mult_B;
  wire       [47:0]   mult_P;
  wire       [7:0]    fixTo_dout;
  wire       [29:0]   tmp_A;
  wire       [17:0]   tmp_B;
  wire       [16:0]   tmp_B_1;
  wire       [5:0]    tmp_shiftRes_1;
  wire       [47:0]   tmp_shiftRes_2;
  wire       [47:0]   tmp_shiftRes_3;
  wire       [47:0]   multRes;
  wire       [47:0]   tmp_shiftRes;
  reg        [47:0]   shiftRes;
  reg        [7:0]    fixTo_dout_regNextWhen;

  assign tmp_A = {{6{din[23]}}, din};
  assign tmp_B_1 = {1'b0,scalerBase};
  assign tmp_B = {{1{tmp_B_1[16]}}, tmp_B_1};
  assign tmp_shiftRes_1 = (scalerExpr - 6'h01);
  assign tmp_shiftRes_2 = ($signed(tmp_shiftRes) + $signed(tmp_shiftRes_3));
  assign tmp_shiftRes_3 = 48'h000000000001;
  AMultB mult (
    .A        (mult_A[29:0]  ), //i
    .B        (mult_B[17:0]  ), //i
    .P        (mult_P[47:0]  ), //o
    .CEs_0    (CEs_0         ), //i
    .CEs_1    (CEs_1         ), //i
    .CEs_2    (CEs_2         ), //i
    .CEs_3    (CEs_3         ), //i
    .clk      (clk           )  //i
  );
  SInt48fixTo7_0_ROUNDTOINF fixTo (
    .din     (shiftRes[47:0]   ), //i
    .dout    (fixTo_dout[7:0]  )  //o
  );
  assign mult_A = tmp_A;
  assign mult_B = tmp_B;
  assign multRes = mult_P;
  assign tmp_shiftRes = ($signed(multRes) >>> scalerExpr);
  assign dout = fixTo_dout_regNextWhen;
  always @(posedge clk) begin
    if(CEs_4) begin
      shiftRes <= (multRes[tmp_shiftRes_1] ? tmp_shiftRes_2 : tmp_shiftRes);
    end
    if(CEs_5) begin
      fixTo_dout_regNextWhen <= fixTo_dout;
    end
  end


endmodule

module EventM2sPipes_8 (
  input               eventIn_valid,
  output              eventIn_ready,
  output              eventOut_valid,
  input               eventOut_ready,
  output              CEs_0,
  output              CEs_1,
  output              CEs_2,
  output              CEs_3,
  output              CEs_4,
  output              CEs_5,
  input               clk,
  input               reset
);

  wire                events_0_valid;
  reg                 events_0_ready;
  wire                events_1_valid;
  reg                 events_1_ready;
  wire                events_2_valid;
  reg                 events_2_ready;
  wire                events_3_valid;
  reg                 events_3_ready;
  wire                events_4_valid;
  reg                 events_4_ready;
  wire                events_5_valid;
  reg                 events_5_ready;
  wire                events_0_m2sPipe_valid;
  wire                events_0_m2sPipe_ready;
  reg                 events_0_rValid;
  wire                when_Stream_l342;
  wire                events_1_m2sPipe_valid;
  wire                events_1_m2sPipe_ready;
  reg                 events_1_rValid;
  wire                when_Stream_l342_1;
  wire                events_2_m2sPipe_valid;
  wire                events_2_m2sPipe_ready;
  reg                 events_2_rValid;
  wire                when_Stream_l342_2;
  wire                events_3_m2sPipe_valid;
  wire                events_3_m2sPipe_ready;
  reg                 events_3_rValid;
  wire                when_Stream_l342_3;
  wire                events_4_m2sPipe_valid;
  wire                events_4_m2sPipe_ready;
  reg                 events_4_rValid;
  wire                when_Stream_l342_4;
  wire                events_5_m2sPipe_valid;
  wire                events_5_m2sPipe_ready;
  reg                 events_5_rValid;
  wire                when_Stream_l342_5;

  assign CEs_0 = events_0_ready;
  assign CEs_1 = events_1_ready;
  assign CEs_2 = events_2_ready;
  assign CEs_3 = events_3_ready;
  assign CEs_4 = events_4_ready;
  assign CEs_5 = events_5_ready;
  assign events_0_valid = eventIn_valid;
  assign eventIn_ready = events_0_ready;
  always @(*) begin
    events_0_ready = events_0_m2sPipe_ready;
    if(when_Stream_l342) begin
      events_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! events_0_m2sPipe_valid);
  assign events_0_m2sPipe_valid = events_0_rValid;
  assign events_1_valid = events_0_m2sPipe_valid;
  assign events_0_m2sPipe_ready = events_1_ready;
  always @(*) begin
    events_1_ready = events_1_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      events_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! events_1_m2sPipe_valid);
  assign events_1_m2sPipe_valid = events_1_rValid;
  assign events_2_valid = events_1_m2sPipe_valid;
  assign events_1_m2sPipe_ready = events_2_ready;
  always @(*) begin
    events_2_ready = events_2_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      events_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! events_2_m2sPipe_valid);
  assign events_2_m2sPipe_valid = events_2_rValid;
  assign events_3_valid = events_2_m2sPipe_valid;
  assign events_2_m2sPipe_ready = events_3_ready;
  always @(*) begin
    events_3_ready = events_3_m2sPipe_ready;
    if(when_Stream_l342_3) begin
      events_3_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! events_3_m2sPipe_valid);
  assign events_3_m2sPipe_valid = events_3_rValid;
  assign events_4_valid = events_3_m2sPipe_valid;
  assign events_3_m2sPipe_ready = events_4_ready;
  always @(*) begin
    events_4_ready = events_4_m2sPipe_ready;
    if(when_Stream_l342_4) begin
      events_4_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! events_4_m2sPipe_valid);
  assign events_4_m2sPipe_valid = events_4_rValid;
  assign events_5_valid = events_4_m2sPipe_valid;
  assign events_4_m2sPipe_ready = events_5_ready;
  always @(*) begin
    events_5_ready = events_5_m2sPipe_ready;
    if(when_Stream_l342_5) begin
      events_5_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! events_5_m2sPipe_valid);
  assign events_5_m2sPipe_valid = events_5_rValid;
  assign eventOut_valid = events_5_m2sPipe_valid;
  assign events_5_m2sPipe_ready = eventOut_ready;
  always @(posedge clk) begin
    if(reset) begin
      events_0_rValid <= 1'b0;
      events_1_rValid <= 1'b0;
      events_2_rValid <= 1'b0;
      events_3_rValid <= 1'b0;
      events_4_rValid <= 1'b0;
      events_5_rValid <= 1'b0;
    end else begin
      if(events_0_ready) begin
        events_0_rValid <= events_0_valid;
      end
      if(events_1_ready) begin
        events_1_rValid <= events_1_valid;
      end
      if(events_2_ready) begin
        events_2_rValid <= events_2_valid;
      end
      if(events_3_ready) begin
        events_3_rValid <= events_3_valid;
      end
      if(events_4_ready) begin
        events_4_rValid <= events_4_valid;
      end
      if(events_5_ready) begin
        events_5_rValid <= events_5_valid;
      end
    end
  end


endmodule

module StreamDemux (
  input      [2:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_0_0_0_0,
  input      [7:0]    io_input_payload_0_0_0_1,
  input      [7:0]    io_input_payload_0_0_0_2,
  input      [7:0]    io_input_payload_0_0_0_3,
  input      [7:0]    io_input_payload_0_0_0_4,
  input      [7:0]    io_input_payload_0_0_0_5,
  input      [7:0]    io_input_payload_0_0_0_6,
  input      [7:0]    io_input_payload_0_0_0_7,
  input      [7:0]    io_input_payload_0_0_0_8,
  input      [7:0]    io_input_payload_0_0_0_9,
  input      [7:0]    io_input_payload_0_0_0_10,
  input      [7:0]    io_input_payload_0_0_0_11,
  input      [7:0]    io_input_payload_0_0_0_12,
  input      [7:0]    io_input_payload_0_0_0_13,
  input      [7:0]    io_input_payload_0_0_0_14,
  input      [7:0]    io_input_payload_0_0_0_15,
  input      [7:0]    io_input_payload_0_0_1_0,
  input      [7:0]    io_input_payload_0_0_1_1,
  input      [7:0]    io_input_payload_0_0_1_2,
  input      [7:0]    io_input_payload_0_0_1_3,
  input      [7:0]    io_input_payload_0_0_1_4,
  input      [7:0]    io_input_payload_0_0_1_5,
  input      [7:0]    io_input_payload_0_0_1_6,
  input      [7:0]    io_input_payload_0_0_1_7,
  input      [7:0]    io_input_payload_0_0_1_8,
  input      [7:0]    io_input_payload_0_0_1_9,
  input      [7:0]    io_input_payload_0_0_1_10,
  input      [7:0]    io_input_payload_0_0_1_11,
  input      [7:0]    io_input_payload_0_0_1_12,
  input      [7:0]    io_input_payload_0_0_1_13,
  input      [7:0]    io_input_payload_0_0_1_14,
  input      [7:0]    io_input_payload_0_0_1_15,
  input      [7:0]    io_input_payload_0_0_2_0,
  input      [7:0]    io_input_payload_0_0_2_1,
  input      [7:0]    io_input_payload_0_0_2_2,
  input      [7:0]    io_input_payload_0_0_2_3,
  input      [7:0]    io_input_payload_0_0_2_4,
  input      [7:0]    io_input_payload_0_0_2_5,
  input      [7:0]    io_input_payload_0_0_2_6,
  input      [7:0]    io_input_payload_0_0_2_7,
  input      [7:0]    io_input_payload_0_0_2_8,
  input      [7:0]    io_input_payload_0_0_2_9,
  input      [7:0]    io_input_payload_0_0_2_10,
  input      [7:0]    io_input_payload_0_0_2_11,
  input      [7:0]    io_input_payload_0_0_2_12,
  input      [7:0]    io_input_payload_0_0_2_13,
  input      [7:0]    io_input_payload_0_0_2_14,
  input      [7:0]    io_input_payload_0_0_2_15,
  input      [7:0]    io_input_payload_0_1_0_0,
  input      [7:0]    io_input_payload_0_1_0_1,
  input      [7:0]    io_input_payload_0_1_0_2,
  input      [7:0]    io_input_payload_0_1_0_3,
  input      [7:0]    io_input_payload_0_1_0_4,
  input      [7:0]    io_input_payload_0_1_0_5,
  input      [7:0]    io_input_payload_0_1_0_6,
  input      [7:0]    io_input_payload_0_1_0_7,
  input      [7:0]    io_input_payload_0_1_0_8,
  input      [7:0]    io_input_payload_0_1_0_9,
  input      [7:0]    io_input_payload_0_1_0_10,
  input      [7:0]    io_input_payload_0_1_0_11,
  input      [7:0]    io_input_payload_0_1_0_12,
  input      [7:0]    io_input_payload_0_1_0_13,
  input      [7:0]    io_input_payload_0_1_0_14,
  input      [7:0]    io_input_payload_0_1_0_15,
  input      [7:0]    io_input_payload_0_1_1_0,
  input      [7:0]    io_input_payload_0_1_1_1,
  input      [7:0]    io_input_payload_0_1_1_2,
  input      [7:0]    io_input_payload_0_1_1_3,
  input      [7:0]    io_input_payload_0_1_1_4,
  input      [7:0]    io_input_payload_0_1_1_5,
  input      [7:0]    io_input_payload_0_1_1_6,
  input      [7:0]    io_input_payload_0_1_1_7,
  input      [7:0]    io_input_payload_0_1_1_8,
  input      [7:0]    io_input_payload_0_1_1_9,
  input      [7:0]    io_input_payload_0_1_1_10,
  input      [7:0]    io_input_payload_0_1_1_11,
  input      [7:0]    io_input_payload_0_1_1_12,
  input      [7:0]    io_input_payload_0_1_1_13,
  input      [7:0]    io_input_payload_0_1_1_14,
  input      [7:0]    io_input_payload_0_1_1_15,
  input      [7:0]    io_input_payload_0_1_2_0,
  input      [7:0]    io_input_payload_0_1_2_1,
  input      [7:0]    io_input_payload_0_1_2_2,
  input      [7:0]    io_input_payload_0_1_2_3,
  input      [7:0]    io_input_payload_0_1_2_4,
  input      [7:0]    io_input_payload_0_1_2_5,
  input      [7:0]    io_input_payload_0_1_2_6,
  input      [7:0]    io_input_payload_0_1_2_7,
  input      [7:0]    io_input_payload_0_1_2_8,
  input      [7:0]    io_input_payload_0_1_2_9,
  input      [7:0]    io_input_payload_0_1_2_10,
  input      [7:0]    io_input_payload_0_1_2_11,
  input      [7:0]    io_input_payload_0_1_2_12,
  input      [7:0]    io_input_payload_0_1_2_13,
  input      [7:0]    io_input_payload_0_1_2_14,
  input      [7:0]    io_input_payload_0_1_2_15,
  input      [7:0]    io_input_payload_0_2_0_0,
  input      [7:0]    io_input_payload_0_2_0_1,
  input      [7:0]    io_input_payload_0_2_0_2,
  input      [7:0]    io_input_payload_0_2_0_3,
  input      [7:0]    io_input_payload_0_2_0_4,
  input      [7:0]    io_input_payload_0_2_0_5,
  input      [7:0]    io_input_payload_0_2_0_6,
  input      [7:0]    io_input_payload_0_2_0_7,
  input      [7:0]    io_input_payload_0_2_0_8,
  input      [7:0]    io_input_payload_0_2_0_9,
  input      [7:0]    io_input_payload_0_2_0_10,
  input      [7:0]    io_input_payload_0_2_0_11,
  input      [7:0]    io_input_payload_0_2_0_12,
  input      [7:0]    io_input_payload_0_2_0_13,
  input      [7:0]    io_input_payload_0_2_0_14,
  input      [7:0]    io_input_payload_0_2_0_15,
  input      [7:0]    io_input_payload_0_2_1_0,
  input      [7:0]    io_input_payload_0_2_1_1,
  input      [7:0]    io_input_payload_0_2_1_2,
  input      [7:0]    io_input_payload_0_2_1_3,
  input      [7:0]    io_input_payload_0_2_1_4,
  input      [7:0]    io_input_payload_0_2_1_5,
  input      [7:0]    io_input_payload_0_2_1_6,
  input      [7:0]    io_input_payload_0_2_1_7,
  input      [7:0]    io_input_payload_0_2_1_8,
  input      [7:0]    io_input_payload_0_2_1_9,
  input      [7:0]    io_input_payload_0_2_1_10,
  input      [7:0]    io_input_payload_0_2_1_11,
  input      [7:0]    io_input_payload_0_2_1_12,
  input      [7:0]    io_input_payload_0_2_1_13,
  input      [7:0]    io_input_payload_0_2_1_14,
  input      [7:0]    io_input_payload_0_2_1_15,
  input      [7:0]    io_input_payload_0_2_2_0,
  input      [7:0]    io_input_payload_0_2_2_1,
  input      [7:0]    io_input_payload_0_2_2_2,
  input      [7:0]    io_input_payload_0_2_2_3,
  input      [7:0]    io_input_payload_0_2_2_4,
  input      [7:0]    io_input_payload_0_2_2_5,
  input      [7:0]    io_input_payload_0_2_2_6,
  input      [7:0]    io_input_payload_0_2_2_7,
  input      [7:0]    io_input_payload_0_2_2_8,
  input      [7:0]    io_input_payload_0_2_2_9,
  input      [7:0]    io_input_payload_0_2_2_10,
  input      [7:0]    io_input_payload_0_2_2_11,
  input      [7:0]    io_input_payload_0_2_2_12,
  input      [7:0]    io_input_payload_0_2_2_13,
  input      [7:0]    io_input_payload_0_2_2_14,
  input      [7:0]    io_input_payload_0_2_2_15,
  input      [7:0]    io_input_payload_1_0_0_0,
  input      [7:0]    io_input_payload_1_0_0_1,
  input      [7:0]    io_input_payload_1_0_0_2,
  input      [7:0]    io_input_payload_1_0_0_3,
  input      [7:0]    io_input_payload_1_0_0_4,
  input      [7:0]    io_input_payload_1_0_0_5,
  input      [7:0]    io_input_payload_1_0_0_6,
  input      [7:0]    io_input_payload_1_0_0_7,
  input      [7:0]    io_input_payload_1_0_0_8,
  input      [7:0]    io_input_payload_1_0_0_9,
  input      [7:0]    io_input_payload_1_0_0_10,
  input      [7:0]    io_input_payload_1_0_0_11,
  input      [7:0]    io_input_payload_1_0_0_12,
  input      [7:0]    io_input_payload_1_0_0_13,
  input      [7:0]    io_input_payload_1_0_0_14,
  input      [7:0]    io_input_payload_1_0_0_15,
  input      [7:0]    io_input_payload_1_0_1_0,
  input      [7:0]    io_input_payload_1_0_1_1,
  input      [7:0]    io_input_payload_1_0_1_2,
  input      [7:0]    io_input_payload_1_0_1_3,
  input      [7:0]    io_input_payload_1_0_1_4,
  input      [7:0]    io_input_payload_1_0_1_5,
  input      [7:0]    io_input_payload_1_0_1_6,
  input      [7:0]    io_input_payload_1_0_1_7,
  input      [7:0]    io_input_payload_1_0_1_8,
  input      [7:0]    io_input_payload_1_0_1_9,
  input      [7:0]    io_input_payload_1_0_1_10,
  input      [7:0]    io_input_payload_1_0_1_11,
  input      [7:0]    io_input_payload_1_0_1_12,
  input      [7:0]    io_input_payload_1_0_1_13,
  input      [7:0]    io_input_payload_1_0_1_14,
  input      [7:0]    io_input_payload_1_0_1_15,
  input      [7:0]    io_input_payload_1_0_2_0,
  input      [7:0]    io_input_payload_1_0_2_1,
  input      [7:0]    io_input_payload_1_0_2_2,
  input      [7:0]    io_input_payload_1_0_2_3,
  input      [7:0]    io_input_payload_1_0_2_4,
  input      [7:0]    io_input_payload_1_0_2_5,
  input      [7:0]    io_input_payload_1_0_2_6,
  input      [7:0]    io_input_payload_1_0_2_7,
  input      [7:0]    io_input_payload_1_0_2_8,
  input      [7:0]    io_input_payload_1_0_2_9,
  input      [7:0]    io_input_payload_1_0_2_10,
  input      [7:0]    io_input_payload_1_0_2_11,
  input      [7:0]    io_input_payload_1_0_2_12,
  input      [7:0]    io_input_payload_1_0_2_13,
  input      [7:0]    io_input_payload_1_0_2_14,
  input      [7:0]    io_input_payload_1_0_2_15,
  input      [7:0]    io_input_payload_1_1_0_0,
  input      [7:0]    io_input_payload_1_1_0_1,
  input      [7:0]    io_input_payload_1_1_0_2,
  input      [7:0]    io_input_payload_1_1_0_3,
  input      [7:0]    io_input_payload_1_1_0_4,
  input      [7:0]    io_input_payload_1_1_0_5,
  input      [7:0]    io_input_payload_1_1_0_6,
  input      [7:0]    io_input_payload_1_1_0_7,
  input      [7:0]    io_input_payload_1_1_0_8,
  input      [7:0]    io_input_payload_1_1_0_9,
  input      [7:0]    io_input_payload_1_1_0_10,
  input      [7:0]    io_input_payload_1_1_0_11,
  input      [7:0]    io_input_payload_1_1_0_12,
  input      [7:0]    io_input_payload_1_1_0_13,
  input      [7:0]    io_input_payload_1_1_0_14,
  input      [7:0]    io_input_payload_1_1_0_15,
  input      [7:0]    io_input_payload_1_1_1_0,
  input      [7:0]    io_input_payload_1_1_1_1,
  input      [7:0]    io_input_payload_1_1_1_2,
  input      [7:0]    io_input_payload_1_1_1_3,
  input      [7:0]    io_input_payload_1_1_1_4,
  input      [7:0]    io_input_payload_1_1_1_5,
  input      [7:0]    io_input_payload_1_1_1_6,
  input      [7:0]    io_input_payload_1_1_1_7,
  input      [7:0]    io_input_payload_1_1_1_8,
  input      [7:0]    io_input_payload_1_1_1_9,
  input      [7:0]    io_input_payload_1_1_1_10,
  input      [7:0]    io_input_payload_1_1_1_11,
  input      [7:0]    io_input_payload_1_1_1_12,
  input      [7:0]    io_input_payload_1_1_1_13,
  input      [7:0]    io_input_payload_1_1_1_14,
  input      [7:0]    io_input_payload_1_1_1_15,
  input      [7:0]    io_input_payload_1_1_2_0,
  input      [7:0]    io_input_payload_1_1_2_1,
  input      [7:0]    io_input_payload_1_1_2_2,
  input      [7:0]    io_input_payload_1_1_2_3,
  input      [7:0]    io_input_payload_1_1_2_4,
  input      [7:0]    io_input_payload_1_1_2_5,
  input      [7:0]    io_input_payload_1_1_2_6,
  input      [7:0]    io_input_payload_1_1_2_7,
  input      [7:0]    io_input_payload_1_1_2_8,
  input      [7:0]    io_input_payload_1_1_2_9,
  input      [7:0]    io_input_payload_1_1_2_10,
  input      [7:0]    io_input_payload_1_1_2_11,
  input      [7:0]    io_input_payload_1_1_2_12,
  input      [7:0]    io_input_payload_1_1_2_13,
  input      [7:0]    io_input_payload_1_1_2_14,
  input      [7:0]    io_input_payload_1_1_2_15,
  input      [7:0]    io_input_payload_1_2_0_0,
  input      [7:0]    io_input_payload_1_2_0_1,
  input      [7:0]    io_input_payload_1_2_0_2,
  input      [7:0]    io_input_payload_1_2_0_3,
  input      [7:0]    io_input_payload_1_2_0_4,
  input      [7:0]    io_input_payload_1_2_0_5,
  input      [7:0]    io_input_payload_1_2_0_6,
  input      [7:0]    io_input_payload_1_2_0_7,
  input      [7:0]    io_input_payload_1_2_0_8,
  input      [7:0]    io_input_payload_1_2_0_9,
  input      [7:0]    io_input_payload_1_2_0_10,
  input      [7:0]    io_input_payload_1_2_0_11,
  input      [7:0]    io_input_payload_1_2_0_12,
  input      [7:0]    io_input_payload_1_2_0_13,
  input      [7:0]    io_input_payload_1_2_0_14,
  input      [7:0]    io_input_payload_1_2_0_15,
  input      [7:0]    io_input_payload_1_2_1_0,
  input      [7:0]    io_input_payload_1_2_1_1,
  input      [7:0]    io_input_payload_1_2_1_2,
  input      [7:0]    io_input_payload_1_2_1_3,
  input      [7:0]    io_input_payload_1_2_1_4,
  input      [7:0]    io_input_payload_1_2_1_5,
  input      [7:0]    io_input_payload_1_2_1_6,
  input      [7:0]    io_input_payload_1_2_1_7,
  input      [7:0]    io_input_payload_1_2_1_8,
  input      [7:0]    io_input_payload_1_2_1_9,
  input      [7:0]    io_input_payload_1_2_1_10,
  input      [7:0]    io_input_payload_1_2_1_11,
  input      [7:0]    io_input_payload_1_2_1_12,
  input      [7:0]    io_input_payload_1_2_1_13,
  input      [7:0]    io_input_payload_1_2_1_14,
  input      [7:0]    io_input_payload_1_2_1_15,
  input      [7:0]    io_input_payload_1_2_2_0,
  input      [7:0]    io_input_payload_1_2_2_1,
  input      [7:0]    io_input_payload_1_2_2_2,
  input      [7:0]    io_input_payload_1_2_2_3,
  input      [7:0]    io_input_payload_1_2_2_4,
  input      [7:0]    io_input_payload_1_2_2_5,
  input      [7:0]    io_input_payload_1_2_2_6,
  input      [7:0]    io_input_payload_1_2_2_7,
  input      [7:0]    io_input_payload_1_2_2_8,
  input      [7:0]    io_input_payload_1_2_2_9,
  input      [7:0]    io_input_payload_1_2_2_10,
  input      [7:0]    io_input_payload_1_2_2_11,
  input      [7:0]    io_input_payload_1_2_2_12,
  input      [7:0]    io_input_payload_1_2_2_13,
  input      [7:0]    io_input_payload_1_2_2_14,
  input      [7:0]    io_input_payload_1_2_2_15,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_0_0_0_0,
  output     [7:0]    io_outputs_0_payload_0_0_0_1,
  output     [7:0]    io_outputs_0_payload_0_0_0_2,
  output     [7:0]    io_outputs_0_payload_0_0_0_3,
  output     [7:0]    io_outputs_0_payload_0_0_0_4,
  output     [7:0]    io_outputs_0_payload_0_0_0_5,
  output     [7:0]    io_outputs_0_payload_0_0_0_6,
  output     [7:0]    io_outputs_0_payload_0_0_0_7,
  output     [7:0]    io_outputs_0_payload_0_0_0_8,
  output     [7:0]    io_outputs_0_payload_0_0_0_9,
  output     [7:0]    io_outputs_0_payload_0_0_0_10,
  output     [7:0]    io_outputs_0_payload_0_0_0_11,
  output     [7:0]    io_outputs_0_payload_0_0_0_12,
  output     [7:0]    io_outputs_0_payload_0_0_0_13,
  output     [7:0]    io_outputs_0_payload_0_0_0_14,
  output     [7:0]    io_outputs_0_payload_0_0_0_15,
  output     [7:0]    io_outputs_0_payload_0_0_1_0,
  output     [7:0]    io_outputs_0_payload_0_0_1_1,
  output     [7:0]    io_outputs_0_payload_0_0_1_2,
  output     [7:0]    io_outputs_0_payload_0_0_1_3,
  output     [7:0]    io_outputs_0_payload_0_0_1_4,
  output     [7:0]    io_outputs_0_payload_0_0_1_5,
  output     [7:0]    io_outputs_0_payload_0_0_1_6,
  output     [7:0]    io_outputs_0_payload_0_0_1_7,
  output     [7:0]    io_outputs_0_payload_0_0_1_8,
  output     [7:0]    io_outputs_0_payload_0_0_1_9,
  output     [7:0]    io_outputs_0_payload_0_0_1_10,
  output     [7:0]    io_outputs_0_payload_0_0_1_11,
  output     [7:0]    io_outputs_0_payload_0_0_1_12,
  output     [7:0]    io_outputs_0_payload_0_0_1_13,
  output     [7:0]    io_outputs_0_payload_0_0_1_14,
  output     [7:0]    io_outputs_0_payload_0_0_1_15,
  output     [7:0]    io_outputs_0_payload_0_0_2_0,
  output     [7:0]    io_outputs_0_payload_0_0_2_1,
  output     [7:0]    io_outputs_0_payload_0_0_2_2,
  output     [7:0]    io_outputs_0_payload_0_0_2_3,
  output     [7:0]    io_outputs_0_payload_0_0_2_4,
  output     [7:0]    io_outputs_0_payload_0_0_2_5,
  output     [7:0]    io_outputs_0_payload_0_0_2_6,
  output     [7:0]    io_outputs_0_payload_0_0_2_7,
  output     [7:0]    io_outputs_0_payload_0_0_2_8,
  output     [7:0]    io_outputs_0_payload_0_0_2_9,
  output     [7:0]    io_outputs_0_payload_0_0_2_10,
  output     [7:0]    io_outputs_0_payload_0_0_2_11,
  output     [7:0]    io_outputs_0_payload_0_0_2_12,
  output     [7:0]    io_outputs_0_payload_0_0_2_13,
  output     [7:0]    io_outputs_0_payload_0_0_2_14,
  output     [7:0]    io_outputs_0_payload_0_0_2_15,
  output     [7:0]    io_outputs_0_payload_0_1_0_0,
  output     [7:0]    io_outputs_0_payload_0_1_0_1,
  output     [7:0]    io_outputs_0_payload_0_1_0_2,
  output     [7:0]    io_outputs_0_payload_0_1_0_3,
  output     [7:0]    io_outputs_0_payload_0_1_0_4,
  output     [7:0]    io_outputs_0_payload_0_1_0_5,
  output     [7:0]    io_outputs_0_payload_0_1_0_6,
  output     [7:0]    io_outputs_0_payload_0_1_0_7,
  output     [7:0]    io_outputs_0_payload_0_1_0_8,
  output     [7:0]    io_outputs_0_payload_0_1_0_9,
  output     [7:0]    io_outputs_0_payload_0_1_0_10,
  output     [7:0]    io_outputs_0_payload_0_1_0_11,
  output     [7:0]    io_outputs_0_payload_0_1_0_12,
  output     [7:0]    io_outputs_0_payload_0_1_0_13,
  output     [7:0]    io_outputs_0_payload_0_1_0_14,
  output     [7:0]    io_outputs_0_payload_0_1_0_15,
  output     [7:0]    io_outputs_0_payload_0_1_1_0,
  output     [7:0]    io_outputs_0_payload_0_1_1_1,
  output     [7:0]    io_outputs_0_payload_0_1_1_2,
  output     [7:0]    io_outputs_0_payload_0_1_1_3,
  output     [7:0]    io_outputs_0_payload_0_1_1_4,
  output     [7:0]    io_outputs_0_payload_0_1_1_5,
  output     [7:0]    io_outputs_0_payload_0_1_1_6,
  output     [7:0]    io_outputs_0_payload_0_1_1_7,
  output     [7:0]    io_outputs_0_payload_0_1_1_8,
  output     [7:0]    io_outputs_0_payload_0_1_1_9,
  output     [7:0]    io_outputs_0_payload_0_1_1_10,
  output     [7:0]    io_outputs_0_payload_0_1_1_11,
  output     [7:0]    io_outputs_0_payload_0_1_1_12,
  output     [7:0]    io_outputs_0_payload_0_1_1_13,
  output     [7:0]    io_outputs_0_payload_0_1_1_14,
  output     [7:0]    io_outputs_0_payload_0_1_1_15,
  output     [7:0]    io_outputs_0_payload_0_1_2_0,
  output     [7:0]    io_outputs_0_payload_0_1_2_1,
  output     [7:0]    io_outputs_0_payload_0_1_2_2,
  output     [7:0]    io_outputs_0_payload_0_1_2_3,
  output     [7:0]    io_outputs_0_payload_0_1_2_4,
  output     [7:0]    io_outputs_0_payload_0_1_2_5,
  output     [7:0]    io_outputs_0_payload_0_1_2_6,
  output     [7:0]    io_outputs_0_payload_0_1_2_7,
  output     [7:0]    io_outputs_0_payload_0_1_2_8,
  output     [7:0]    io_outputs_0_payload_0_1_2_9,
  output     [7:0]    io_outputs_0_payload_0_1_2_10,
  output     [7:0]    io_outputs_0_payload_0_1_2_11,
  output     [7:0]    io_outputs_0_payload_0_1_2_12,
  output     [7:0]    io_outputs_0_payload_0_1_2_13,
  output     [7:0]    io_outputs_0_payload_0_1_2_14,
  output     [7:0]    io_outputs_0_payload_0_1_2_15,
  output     [7:0]    io_outputs_0_payload_0_2_0_0,
  output     [7:0]    io_outputs_0_payload_0_2_0_1,
  output     [7:0]    io_outputs_0_payload_0_2_0_2,
  output     [7:0]    io_outputs_0_payload_0_2_0_3,
  output     [7:0]    io_outputs_0_payload_0_2_0_4,
  output     [7:0]    io_outputs_0_payload_0_2_0_5,
  output     [7:0]    io_outputs_0_payload_0_2_0_6,
  output     [7:0]    io_outputs_0_payload_0_2_0_7,
  output     [7:0]    io_outputs_0_payload_0_2_0_8,
  output     [7:0]    io_outputs_0_payload_0_2_0_9,
  output     [7:0]    io_outputs_0_payload_0_2_0_10,
  output     [7:0]    io_outputs_0_payload_0_2_0_11,
  output     [7:0]    io_outputs_0_payload_0_2_0_12,
  output     [7:0]    io_outputs_0_payload_0_2_0_13,
  output     [7:0]    io_outputs_0_payload_0_2_0_14,
  output     [7:0]    io_outputs_0_payload_0_2_0_15,
  output     [7:0]    io_outputs_0_payload_0_2_1_0,
  output     [7:0]    io_outputs_0_payload_0_2_1_1,
  output     [7:0]    io_outputs_0_payload_0_2_1_2,
  output     [7:0]    io_outputs_0_payload_0_2_1_3,
  output     [7:0]    io_outputs_0_payload_0_2_1_4,
  output     [7:0]    io_outputs_0_payload_0_2_1_5,
  output     [7:0]    io_outputs_0_payload_0_2_1_6,
  output     [7:0]    io_outputs_0_payload_0_2_1_7,
  output     [7:0]    io_outputs_0_payload_0_2_1_8,
  output     [7:0]    io_outputs_0_payload_0_2_1_9,
  output     [7:0]    io_outputs_0_payload_0_2_1_10,
  output     [7:0]    io_outputs_0_payload_0_2_1_11,
  output     [7:0]    io_outputs_0_payload_0_2_1_12,
  output     [7:0]    io_outputs_0_payload_0_2_1_13,
  output     [7:0]    io_outputs_0_payload_0_2_1_14,
  output     [7:0]    io_outputs_0_payload_0_2_1_15,
  output     [7:0]    io_outputs_0_payload_0_2_2_0,
  output     [7:0]    io_outputs_0_payload_0_2_2_1,
  output     [7:0]    io_outputs_0_payload_0_2_2_2,
  output     [7:0]    io_outputs_0_payload_0_2_2_3,
  output     [7:0]    io_outputs_0_payload_0_2_2_4,
  output     [7:0]    io_outputs_0_payload_0_2_2_5,
  output     [7:0]    io_outputs_0_payload_0_2_2_6,
  output     [7:0]    io_outputs_0_payload_0_2_2_7,
  output     [7:0]    io_outputs_0_payload_0_2_2_8,
  output     [7:0]    io_outputs_0_payload_0_2_2_9,
  output     [7:0]    io_outputs_0_payload_0_2_2_10,
  output     [7:0]    io_outputs_0_payload_0_2_2_11,
  output     [7:0]    io_outputs_0_payload_0_2_2_12,
  output     [7:0]    io_outputs_0_payload_0_2_2_13,
  output     [7:0]    io_outputs_0_payload_0_2_2_14,
  output     [7:0]    io_outputs_0_payload_0_2_2_15,
  output     [7:0]    io_outputs_0_payload_1_0_0_0,
  output     [7:0]    io_outputs_0_payload_1_0_0_1,
  output     [7:0]    io_outputs_0_payload_1_0_0_2,
  output     [7:0]    io_outputs_0_payload_1_0_0_3,
  output     [7:0]    io_outputs_0_payload_1_0_0_4,
  output     [7:0]    io_outputs_0_payload_1_0_0_5,
  output     [7:0]    io_outputs_0_payload_1_0_0_6,
  output     [7:0]    io_outputs_0_payload_1_0_0_7,
  output     [7:0]    io_outputs_0_payload_1_0_0_8,
  output     [7:0]    io_outputs_0_payload_1_0_0_9,
  output     [7:0]    io_outputs_0_payload_1_0_0_10,
  output     [7:0]    io_outputs_0_payload_1_0_0_11,
  output     [7:0]    io_outputs_0_payload_1_0_0_12,
  output     [7:0]    io_outputs_0_payload_1_0_0_13,
  output     [7:0]    io_outputs_0_payload_1_0_0_14,
  output     [7:0]    io_outputs_0_payload_1_0_0_15,
  output     [7:0]    io_outputs_0_payload_1_0_1_0,
  output     [7:0]    io_outputs_0_payload_1_0_1_1,
  output     [7:0]    io_outputs_0_payload_1_0_1_2,
  output     [7:0]    io_outputs_0_payload_1_0_1_3,
  output     [7:0]    io_outputs_0_payload_1_0_1_4,
  output     [7:0]    io_outputs_0_payload_1_0_1_5,
  output     [7:0]    io_outputs_0_payload_1_0_1_6,
  output     [7:0]    io_outputs_0_payload_1_0_1_7,
  output     [7:0]    io_outputs_0_payload_1_0_1_8,
  output     [7:0]    io_outputs_0_payload_1_0_1_9,
  output     [7:0]    io_outputs_0_payload_1_0_1_10,
  output     [7:0]    io_outputs_0_payload_1_0_1_11,
  output     [7:0]    io_outputs_0_payload_1_0_1_12,
  output     [7:0]    io_outputs_0_payload_1_0_1_13,
  output     [7:0]    io_outputs_0_payload_1_0_1_14,
  output     [7:0]    io_outputs_0_payload_1_0_1_15,
  output     [7:0]    io_outputs_0_payload_1_0_2_0,
  output     [7:0]    io_outputs_0_payload_1_0_2_1,
  output     [7:0]    io_outputs_0_payload_1_0_2_2,
  output     [7:0]    io_outputs_0_payload_1_0_2_3,
  output     [7:0]    io_outputs_0_payload_1_0_2_4,
  output     [7:0]    io_outputs_0_payload_1_0_2_5,
  output     [7:0]    io_outputs_0_payload_1_0_2_6,
  output     [7:0]    io_outputs_0_payload_1_0_2_7,
  output     [7:0]    io_outputs_0_payload_1_0_2_8,
  output     [7:0]    io_outputs_0_payload_1_0_2_9,
  output     [7:0]    io_outputs_0_payload_1_0_2_10,
  output     [7:0]    io_outputs_0_payload_1_0_2_11,
  output     [7:0]    io_outputs_0_payload_1_0_2_12,
  output     [7:0]    io_outputs_0_payload_1_0_2_13,
  output     [7:0]    io_outputs_0_payload_1_0_2_14,
  output     [7:0]    io_outputs_0_payload_1_0_2_15,
  output     [7:0]    io_outputs_0_payload_1_1_0_0,
  output     [7:0]    io_outputs_0_payload_1_1_0_1,
  output     [7:0]    io_outputs_0_payload_1_1_0_2,
  output     [7:0]    io_outputs_0_payload_1_1_0_3,
  output     [7:0]    io_outputs_0_payload_1_1_0_4,
  output     [7:0]    io_outputs_0_payload_1_1_0_5,
  output     [7:0]    io_outputs_0_payload_1_1_0_6,
  output     [7:0]    io_outputs_0_payload_1_1_0_7,
  output     [7:0]    io_outputs_0_payload_1_1_0_8,
  output     [7:0]    io_outputs_0_payload_1_1_0_9,
  output     [7:0]    io_outputs_0_payload_1_1_0_10,
  output     [7:0]    io_outputs_0_payload_1_1_0_11,
  output     [7:0]    io_outputs_0_payload_1_1_0_12,
  output     [7:0]    io_outputs_0_payload_1_1_0_13,
  output     [7:0]    io_outputs_0_payload_1_1_0_14,
  output     [7:0]    io_outputs_0_payload_1_1_0_15,
  output     [7:0]    io_outputs_0_payload_1_1_1_0,
  output     [7:0]    io_outputs_0_payload_1_1_1_1,
  output     [7:0]    io_outputs_0_payload_1_1_1_2,
  output     [7:0]    io_outputs_0_payload_1_1_1_3,
  output     [7:0]    io_outputs_0_payload_1_1_1_4,
  output     [7:0]    io_outputs_0_payload_1_1_1_5,
  output     [7:0]    io_outputs_0_payload_1_1_1_6,
  output     [7:0]    io_outputs_0_payload_1_1_1_7,
  output     [7:0]    io_outputs_0_payload_1_1_1_8,
  output     [7:0]    io_outputs_0_payload_1_1_1_9,
  output     [7:0]    io_outputs_0_payload_1_1_1_10,
  output     [7:0]    io_outputs_0_payload_1_1_1_11,
  output     [7:0]    io_outputs_0_payload_1_1_1_12,
  output     [7:0]    io_outputs_0_payload_1_1_1_13,
  output     [7:0]    io_outputs_0_payload_1_1_1_14,
  output     [7:0]    io_outputs_0_payload_1_1_1_15,
  output     [7:0]    io_outputs_0_payload_1_1_2_0,
  output     [7:0]    io_outputs_0_payload_1_1_2_1,
  output     [7:0]    io_outputs_0_payload_1_1_2_2,
  output     [7:0]    io_outputs_0_payload_1_1_2_3,
  output     [7:0]    io_outputs_0_payload_1_1_2_4,
  output     [7:0]    io_outputs_0_payload_1_1_2_5,
  output     [7:0]    io_outputs_0_payload_1_1_2_6,
  output     [7:0]    io_outputs_0_payload_1_1_2_7,
  output     [7:0]    io_outputs_0_payload_1_1_2_8,
  output     [7:0]    io_outputs_0_payload_1_1_2_9,
  output     [7:0]    io_outputs_0_payload_1_1_2_10,
  output     [7:0]    io_outputs_0_payload_1_1_2_11,
  output     [7:0]    io_outputs_0_payload_1_1_2_12,
  output     [7:0]    io_outputs_0_payload_1_1_2_13,
  output     [7:0]    io_outputs_0_payload_1_1_2_14,
  output     [7:0]    io_outputs_0_payload_1_1_2_15,
  output     [7:0]    io_outputs_0_payload_1_2_0_0,
  output     [7:0]    io_outputs_0_payload_1_2_0_1,
  output     [7:0]    io_outputs_0_payload_1_2_0_2,
  output     [7:0]    io_outputs_0_payload_1_2_0_3,
  output     [7:0]    io_outputs_0_payload_1_2_0_4,
  output     [7:0]    io_outputs_0_payload_1_2_0_5,
  output     [7:0]    io_outputs_0_payload_1_2_0_6,
  output     [7:0]    io_outputs_0_payload_1_2_0_7,
  output     [7:0]    io_outputs_0_payload_1_2_0_8,
  output     [7:0]    io_outputs_0_payload_1_2_0_9,
  output     [7:0]    io_outputs_0_payload_1_2_0_10,
  output     [7:0]    io_outputs_0_payload_1_2_0_11,
  output     [7:0]    io_outputs_0_payload_1_2_0_12,
  output     [7:0]    io_outputs_0_payload_1_2_0_13,
  output     [7:0]    io_outputs_0_payload_1_2_0_14,
  output     [7:0]    io_outputs_0_payload_1_2_0_15,
  output     [7:0]    io_outputs_0_payload_1_2_1_0,
  output     [7:0]    io_outputs_0_payload_1_2_1_1,
  output     [7:0]    io_outputs_0_payload_1_2_1_2,
  output     [7:0]    io_outputs_0_payload_1_2_1_3,
  output     [7:0]    io_outputs_0_payload_1_2_1_4,
  output     [7:0]    io_outputs_0_payload_1_2_1_5,
  output     [7:0]    io_outputs_0_payload_1_2_1_6,
  output     [7:0]    io_outputs_0_payload_1_2_1_7,
  output     [7:0]    io_outputs_0_payload_1_2_1_8,
  output     [7:0]    io_outputs_0_payload_1_2_1_9,
  output     [7:0]    io_outputs_0_payload_1_2_1_10,
  output     [7:0]    io_outputs_0_payload_1_2_1_11,
  output     [7:0]    io_outputs_0_payload_1_2_1_12,
  output     [7:0]    io_outputs_0_payload_1_2_1_13,
  output     [7:0]    io_outputs_0_payload_1_2_1_14,
  output     [7:0]    io_outputs_0_payload_1_2_1_15,
  output     [7:0]    io_outputs_0_payload_1_2_2_0,
  output     [7:0]    io_outputs_0_payload_1_2_2_1,
  output     [7:0]    io_outputs_0_payload_1_2_2_2,
  output     [7:0]    io_outputs_0_payload_1_2_2_3,
  output     [7:0]    io_outputs_0_payload_1_2_2_4,
  output     [7:0]    io_outputs_0_payload_1_2_2_5,
  output     [7:0]    io_outputs_0_payload_1_2_2_6,
  output     [7:0]    io_outputs_0_payload_1_2_2_7,
  output     [7:0]    io_outputs_0_payload_1_2_2_8,
  output     [7:0]    io_outputs_0_payload_1_2_2_9,
  output     [7:0]    io_outputs_0_payload_1_2_2_10,
  output     [7:0]    io_outputs_0_payload_1_2_2_11,
  output     [7:0]    io_outputs_0_payload_1_2_2_12,
  output     [7:0]    io_outputs_0_payload_1_2_2_13,
  output     [7:0]    io_outputs_0_payload_1_2_2_14,
  output     [7:0]    io_outputs_0_payload_1_2_2_15,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_0_0_0_0,
  output     [7:0]    io_outputs_1_payload_0_0_0_1,
  output     [7:0]    io_outputs_1_payload_0_0_0_2,
  output     [7:0]    io_outputs_1_payload_0_0_0_3,
  output     [7:0]    io_outputs_1_payload_0_0_0_4,
  output     [7:0]    io_outputs_1_payload_0_0_0_5,
  output     [7:0]    io_outputs_1_payload_0_0_0_6,
  output     [7:0]    io_outputs_1_payload_0_0_0_7,
  output     [7:0]    io_outputs_1_payload_0_0_0_8,
  output     [7:0]    io_outputs_1_payload_0_0_0_9,
  output     [7:0]    io_outputs_1_payload_0_0_0_10,
  output     [7:0]    io_outputs_1_payload_0_0_0_11,
  output     [7:0]    io_outputs_1_payload_0_0_0_12,
  output     [7:0]    io_outputs_1_payload_0_0_0_13,
  output     [7:0]    io_outputs_1_payload_0_0_0_14,
  output     [7:0]    io_outputs_1_payload_0_0_0_15,
  output     [7:0]    io_outputs_1_payload_0_0_1_0,
  output     [7:0]    io_outputs_1_payload_0_0_1_1,
  output     [7:0]    io_outputs_1_payload_0_0_1_2,
  output     [7:0]    io_outputs_1_payload_0_0_1_3,
  output     [7:0]    io_outputs_1_payload_0_0_1_4,
  output     [7:0]    io_outputs_1_payload_0_0_1_5,
  output     [7:0]    io_outputs_1_payload_0_0_1_6,
  output     [7:0]    io_outputs_1_payload_0_0_1_7,
  output     [7:0]    io_outputs_1_payload_0_0_1_8,
  output     [7:0]    io_outputs_1_payload_0_0_1_9,
  output     [7:0]    io_outputs_1_payload_0_0_1_10,
  output     [7:0]    io_outputs_1_payload_0_0_1_11,
  output     [7:0]    io_outputs_1_payload_0_0_1_12,
  output     [7:0]    io_outputs_1_payload_0_0_1_13,
  output     [7:0]    io_outputs_1_payload_0_0_1_14,
  output     [7:0]    io_outputs_1_payload_0_0_1_15,
  output     [7:0]    io_outputs_1_payload_0_0_2_0,
  output     [7:0]    io_outputs_1_payload_0_0_2_1,
  output     [7:0]    io_outputs_1_payload_0_0_2_2,
  output     [7:0]    io_outputs_1_payload_0_0_2_3,
  output     [7:0]    io_outputs_1_payload_0_0_2_4,
  output     [7:0]    io_outputs_1_payload_0_0_2_5,
  output     [7:0]    io_outputs_1_payload_0_0_2_6,
  output     [7:0]    io_outputs_1_payload_0_0_2_7,
  output     [7:0]    io_outputs_1_payload_0_0_2_8,
  output     [7:0]    io_outputs_1_payload_0_0_2_9,
  output     [7:0]    io_outputs_1_payload_0_0_2_10,
  output     [7:0]    io_outputs_1_payload_0_0_2_11,
  output     [7:0]    io_outputs_1_payload_0_0_2_12,
  output     [7:0]    io_outputs_1_payload_0_0_2_13,
  output     [7:0]    io_outputs_1_payload_0_0_2_14,
  output     [7:0]    io_outputs_1_payload_0_0_2_15,
  output     [7:0]    io_outputs_1_payload_0_1_0_0,
  output     [7:0]    io_outputs_1_payload_0_1_0_1,
  output     [7:0]    io_outputs_1_payload_0_1_0_2,
  output     [7:0]    io_outputs_1_payload_0_1_0_3,
  output     [7:0]    io_outputs_1_payload_0_1_0_4,
  output     [7:0]    io_outputs_1_payload_0_1_0_5,
  output     [7:0]    io_outputs_1_payload_0_1_0_6,
  output     [7:0]    io_outputs_1_payload_0_1_0_7,
  output     [7:0]    io_outputs_1_payload_0_1_0_8,
  output     [7:0]    io_outputs_1_payload_0_1_0_9,
  output     [7:0]    io_outputs_1_payload_0_1_0_10,
  output     [7:0]    io_outputs_1_payload_0_1_0_11,
  output     [7:0]    io_outputs_1_payload_0_1_0_12,
  output     [7:0]    io_outputs_1_payload_0_1_0_13,
  output     [7:0]    io_outputs_1_payload_0_1_0_14,
  output     [7:0]    io_outputs_1_payload_0_1_0_15,
  output     [7:0]    io_outputs_1_payload_0_1_1_0,
  output     [7:0]    io_outputs_1_payload_0_1_1_1,
  output     [7:0]    io_outputs_1_payload_0_1_1_2,
  output     [7:0]    io_outputs_1_payload_0_1_1_3,
  output     [7:0]    io_outputs_1_payload_0_1_1_4,
  output     [7:0]    io_outputs_1_payload_0_1_1_5,
  output     [7:0]    io_outputs_1_payload_0_1_1_6,
  output     [7:0]    io_outputs_1_payload_0_1_1_7,
  output     [7:0]    io_outputs_1_payload_0_1_1_8,
  output     [7:0]    io_outputs_1_payload_0_1_1_9,
  output     [7:0]    io_outputs_1_payload_0_1_1_10,
  output     [7:0]    io_outputs_1_payload_0_1_1_11,
  output     [7:0]    io_outputs_1_payload_0_1_1_12,
  output     [7:0]    io_outputs_1_payload_0_1_1_13,
  output     [7:0]    io_outputs_1_payload_0_1_1_14,
  output     [7:0]    io_outputs_1_payload_0_1_1_15,
  output     [7:0]    io_outputs_1_payload_0_1_2_0,
  output     [7:0]    io_outputs_1_payload_0_1_2_1,
  output     [7:0]    io_outputs_1_payload_0_1_2_2,
  output     [7:0]    io_outputs_1_payload_0_1_2_3,
  output     [7:0]    io_outputs_1_payload_0_1_2_4,
  output     [7:0]    io_outputs_1_payload_0_1_2_5,
  output     [7:0]    io_outputs_1_payload_0_1_2_6,
  output     [7:0]    io_outputs_1_payload_0_1_2_7,
  output     [7:0]    io_outputs_1_payload_0_1_2_8,
  output     [7:0]    io_outputs_1_payload_0_1_2_9,
  output     [7:0]    io_outputs_1_payload_0_1_2_10,
  output     [7:0]    io_outputs_1_payload_0_1_2_11,
  output     [7:0]    io_outputs_1_payload_0_1_2_12,
  output     [7:0]    io_outputs_1_payload_0_1_2_13,
  output     [7:0]    io_outputs_1_payload_0_1_2_14,
  output     [7:0]    io_outputs_1_payload_0_1_2_15,
  output     [7:0]    io_outputs_1_payload_0_2_0_0,
  output     [7:0]    io_outputs_1_payload_0_2_0_1,
  output     [7:0]    io_outputs_1_payload_0_2_0_2,
  output     [7:0]    io_outputs_1_payload_0_2_0_3,
  output     [7:0]    io_outputs_1_payload_0_2_0_4,
  output     [7:0]    io_outputs_1_payload_0_2_0_5,
  output     [7:0]    io_outputs_1_payload_0_2_0_6,
  output     [7:0]    io_outputs_1_payload_0_2_0_7,
  output     [7:0]    io_outputs_1_payload_0_2_0_8,
  output     [7:0]    io_outputs_1_payload_0_2_0_9,
  output     [7:0]    io_outputs_1_payload_0_2_0_10,
  output     [7:0]    io_outputs_1_payload_0_2_0_11,
  output     [7:0]    io_outputs_1_payload_0_2_0_12,
  output     [7:0]    io_outputs_1_payload_0_2_0_13,
  output     [7:0]    io_outputs_1_payload_0_2_0_14,
  output     [7:0]    io_outputs_1_payload_0_2_0_15,
  output     [7:0]    io_outputs_1_payload_0_2_1_0,
  output     [7:0]    io_outputs_1_payload_0_2_1_1,
  output     [7:0]    io_outputs_1_payload_0_2_1_2,
  output     [7:0]    io_outputs_1_payload_0_2_1_3,
  output     [7:0]    io_outputs_1_payload_0_2_1_4,
  output     [7:0]    io_outputs_1_payload_0_2_1_5,
  output     [7:0]    io_outputs_1_payload_0_2_1_6,
  output     [7:0]    io_outputs_1_payload_0_2_1_7,
  output     [7:0]    io_outputs_1_payload_0_2_1_8,
  output     [7:0]    io_outputs_1_payload_0_2_1_9,
  output     [7:0]    io_outputs_1_payload_0_2_1_10,
  output     [7:0]    io_outputs_1_payload_0_2_1_11,
  output     [7:0]    io_outputs_1_payload_0_2_1_12,
  output     [7:0]    io_outputs_1_payload_0_2_1_13,
  output     [7:0]    io_outputs_1_payload_0_2_1_14,
  output     [7:0]    io_outputs_1_payload_0_2_1_15,
  output     [7:0]    io_outputs_1_payload_0_2_2_0,
  output     [7:0]    io_outputs_1_payload_0_2_2_1,
  output     [7:0]    io_outputs_1_payload_0_2_2_2,
  output     [7:0]    io_outputs_1_payload_0_2_2_3,
  output     [7:0]    io_outputs_1_payload_0_2_2_4,
  output     [7:0]    io_outputs_1_payload_0_2_2_5,
  output     [7:0]    io_outputs_1_payload_0_2_2_6,
  output     [7:0]    io_outputs_1_payload_0_2_2_7,
  output     [7:0]    io_outputs_1_payload_0_2_2_8,
  output     [7:0]    io_outputs_1_payload_0_2_2_9,
  output     [7:0]    io_outputs_1_payload_0_2_2_10,
  output     [7:0]    io_outputs_1_payload_0_2_2_11,
  output     [7:0]    io_outputs_1_payload_0_2_2_12,
  output     [7:0]    io_outputs_1_payload_0_2_2_13,
  output     [7:0]    io_outputs_1_payload_0_2_2_14,
  output     [7:0]    io_outputs_1_payload_0_2_2_15,
  output     [7:0]    io_outputs_1_payload_1_0_0_0,
  output     [7:0]    io_outputs_1_payload_1_0_0_1,
  output     [7:0]    io_outputs_1_payload_1_0_0_2,
  output     [7:0]    io_outputs_1_payload_1_0_0_3,
  output     [7:0]    io_outputs_1_payload_1_0_0_4,
  output     [7:0]    io_outputs_1_payload_1_0_0_5,
  output     [7:0]    io_outputs_1_payload_1_0_0_6,
  output     [7:0]    io_outputs_1_payload_1_0_0_7,
  output     [7:0]    io_outputs_1_payload_1_0_0_8,
  output     [7:0]    io_outputs_1_payload_1_0_0_9,
  output     [7:0]    io_outputs_1_payload_1_0_0_10,
  output     [7:0]    io_outputs_1_payload_1_0_0_11,
  output     [7:0]    io_outputs_1_payload_1_0_0_12,
  output     [7:0]    io_outputs_1_payload_1_0_0_13,
  output     [7:0]    io_outputs_1_payload_1_0_0_14,
  output     [7:0]    io_outputs_1_payload_1_0_0_15,
  output     [7:0]    io_outputs_1_payload_1_0_1_0,
  output     [7:0]    io_outputs_1_payload_1_0_1_1,
  output     [7:0]    io_outputs_1_payload_1_0_1_2,
  output     [7:0]    io_outputs_1_payload_1_0_1_3,
  output     [7:0]    io_outputs_1_payload_1_0_1_4,
  output     [7:0]    io_outputs_1_payload_1_0_1_5,
  output     [7:0]    io_outputs_1_payload_1_0_1_6,
  output     [7:0]    io_outputs_1_payload_1_0_1_7,
  output     [7:0]    io_outputs_1_payload_1_0_1_8,
  output     [7:0]    io_outputs_1_payload_1_0_1_9,
  output     [7:0]    io_outputs_1_payload_1_0_1_10,
  output     [7:0]    io_outputs_1_payload_1_0_1_11,
  output     [7:0]    io_outputs_1_payload_1_0_1_12,
  output     [7:0]    io_outputs_1_payload_1_0_1_13,
  output     [7:0]    io_outputs_1_payload_1_0_1_14,
  output     [7:0]    io_outputs_1_payload_1_0_1_15,
  output     [7:0]    io_outputs_1_payload_1_0_2_0,
  output     [7:0]    io_outputs_1_payload_1_0_2_1,
  output     [7:0]    io_outputs_1_payload_1_0_2_2,
  output     [7:0]    io_outputs_1_payload_1_0_2_3,
  output     [7:0]    io_outputs_1_payload_1_0_2_4,
  output     [7:0]    io_outputs_1_payload_1_0_2_5,
  output     [7:0]    io_outputs_1_payload_1_0_2_6,
  output     [7:0]    io_outputs_1_payload_1_0_2_7,
  output     [7:0]    io_outputs_1_payload_1_0_2_8,
  output     [7:0]    io_outputs_1_payload_1_0_2_9,
  output     [7:0]    io_outputs_1_payload_1_0_2_10,
  output     [7:0]    io_outputs_1_payload_1_0_2_11,
  output     [7:0]    io_outputs_1_payload_1_0_2_12,
  output     [7:0]    io_outputs_1_payload_1_0_2_13,
  output     [7:0]    io_outputs_1_payload_1_0_2_14,
  output     [7:0]    io_outputs_1_payload_1_0_2_15,
  output     [7:0]    io_outputs_1_payload_1_1_0_0,
  output     [7:0]    io_outputs_1_payload_1_1_0_1,
  output     [7:0]    io_outputs_1_payload_1_1_0_2,
  output     [7:0]    io_outputs_1_payload_1_1_0_3,
  output     [7:0]    io_outputs_1_payload_1_1_0_4,
  output     [7:0]    io_outputs_1_payload_1_1_0_5,
  output     [7:0]    io_outputs_1_payload_1_1_0_6,
  output     [7:0]    io_outputs_1_payload_1_1_0_7,
  output     [7:0]    io_outputs_1_payload_1_1_0_8,
  output     [7:0]    io_outputs_1_payload_1_1_0_9,
  output     [7:0]    io_outputs_1_payload_1_1_0_10,
  output     [7:0]    io_outputs_1_payload_1_1_0_11,
  output     [7:0]    io_outputs_1_payload_1_1_0_12,
  output     [7:0]    io_outputs_1_payload_1_1_0_13,
  output     [7:0]    io_outputs_1_payload_1_1_0_14,
  output     [7:0]    io_outputs_1_payload_1_1_0_15,
  output     [7:0]    io_outputs_1_payload_1_1_1_0,
  output     [7:0]    io_outputs_1_payload_1_1_1_1,
  output     [7:0]    io_outputs_1_payload_1_1_1_2,
  output     [7:0]    io_outputs_1_payload_1_1_1_3,
  output     [7:0]    io_outputs_1_payload_1_1_1_4,
  output     [7:0]    io_outputs_1_payload_1_1_1_5,
  output     [7:0]    io_outputs_1_payload_1_1_1_6,
  output     [7:0]    io_outputs_1_payload_1_1_1_7,
  output     [7:0]    io_outputs_1_payload_1_1_1_8,
  output     [7:0]    io_outputs_1_payload_1_1_1_9,
  output     [7:0]    io_outputs_1_payload_1_1_1_10,
  output     [7:0]    io_outputs_1_payload_1_1_1_11,
  output     [7:0]    io_outputs_1_payload_1_1_1_12,
  output     [7:0]    io_outputs_1_payload_1_1_1_13,
  output     [7:0]    io_outputs_1_payload_1_1_1_14,
  output     [7:0]    io_outputs_1_payload_1_1_1_15,
  output     [7:0]    io_outputs_1_payload_1_1_2_0,
  output     [7:0]    io_outputs_1_payload_1_1_2_1,
  output     [7:0]    io_outputs_1_payload_1_1_2_2,
  output     [7:0]    io_outputs_1_payload_1_1_2_3,
  output     [7:0]    io_outputs_1_payload_1_1_2_4,
  output     [7:0]    io_outputs_1_payload_1_1_2_5,
  output     [7:0]    io_outputs_1_payload_1_1_2_6,
  output     [7:0]    io_outputs_1_payload_1_1_2_7,
  output     [7:0]    io_outputs_1_payload_1_1_2_8,
  output     [7:0]    io_outputs_1_payload_1_1_2_9,
  output     [7:0]    io_outputs_1_payload_1_1_2_10,
  output     [7:0]    io_outputs_1_payload_1_1_2_11,
  output     [7:0]    io_outputs_1_payload_1_1_2_12,
  output     [7:0]    io_outputs_1_payload_1_1_2_13,
  output     [7:0]    io_outputs_1_payload_1_1_2_14,
  output     [7:0]    io_outputs_1_payload_1_1_2_15,
  output     [7:0]    io_outputs_1_payload_1_2_0_0,
  output     [7:0]    io_outputs_1_payload_1_2_0_1,
  output     [7:0]    io_outputs_1_payload_1_2_0_2,
  output     [7:0]    io_outputs_1_payload_1_2_0_3,
  output     [7:0]    io_outputs_1_payload_1_2_0_4,
  output     [7:0]    io_outputs_1_payload_1_2_0_5,
  output     [7:0]    io_outputs_1_payload_1_2_0_6,
  output     [7:0]    io_outputs_1_payload_1_2_0_7,
  output     [7:0]    io_outputs_1_payload_1_2_0_8,
  output     [7:0]    io_outputs_1_payload_1_2_0_9,
  output     [7:0]    io_outputs_1_payload_1_2_0_10,
  output     [7:0]    io_outputs_1_payload_1_2_0_11,
  output     [7:0]    io_outputs_1_payload_1_2_0_12,
  output     [7:0]    io_outputs_1_payload_1_2_0_13,
  output     [7:0]    io_outputs_1_payload_1_2_0_14,
  output     [7:0]    io_outputs_1_payload_1_2_0_15,
  output     [7:0]    io_outputs_1_payload_1_2_1_0,
  output     [7:0]    io_outputs_1_payload_1_2_1_1,
  output     [7:0]    io_outputs_1_payload_1_2_1_2,
  output     [7:0]    io_outputs_1_payload_1_2_1_3,
  output     [7:0]    io_outputs_1_payload_1_2_1_4,
  output     [7:0]    io_outputs_1_payload_1_2_1_5,
  output     [7:0]    io_outputs_1_payload_1_2_1_6,
  output     [7:0]    io_outputs_1_payload_1_2_1_7,
  output     [7:0]    io_outputs_1_payload_1_2_1_8,
  output     [7:0]    io_outputs_1_payload_1_2_1_9,
  output     [7:0]    io_outputs_1_payload_1_2_1_10,
  output     [7:0]    io_outputs_1_payload_1_2_1_11,
  output     [7:0]    io_outputs_1_payload_1_2_1_12,
  output     [7:0]    io_outputs_1_payload_1_2_1_13,
  output     [7:0]    io_outputs_1_payload_1_2_1_14,
  output     [7:0]    io_outputs_1_payload_1_2_1_15,
  output     [7:0]    io_outputs_1_payload_1_2_2_0,
  output     [7:0]    io_outputs_1_payload_1_2_2_1,
  output     [7:0]    io_outputs_1_payload_1_2_2_2,
  output     [7:0]    io_outputs_1_payload_1_2_2_3,
  output     [7:0]    io_outputs_1_payload_1_2_2_4,
  output     [7:0]    io_outputs_1_payload_1_2_2_5,
  output     [7:0]    io_outputs_1_payload_1_2_2_6,
  output     [7:0]    io_outputs_1_payload_1_2_2_7,
  output     [7:0]    io_outputs_1_payload_1_2_2_8,
  output     [7:0]    io_outputs_1_payload_1_2_2_9,
  output     [7:0]    io_outputs_1_payload_1_2_2_10,
  output     [7:0]    io_outputs_1_payload_1_2_2_11,
  output     [7:0]    io_outputs_1_payload_1_2_2_12,
  output     [7:0]    io_outputs_1_payload_1_2_2_13,
  output     [7:0]    io_outputs_1_payload_1_2_2_14,
  output     [7:0]    io_outputs_1_payload_1_2_2_15,
  output reg          io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [7:0]    io_outputs_2_payload_0_0_0_0,
  output     [7:0]    io_outputs_2_payload_0_0_0_1,
  output     [7:0]    io_outputs_2_payload_0_0_0_2,
  output     [7:0]    io_outputs_2_payload_0_0_0_3,
  output     [7:0]    io_outputs_2_payload_0_0_0_4,
  output     [7:0]    io_outputs_2_payload_0_0_0_5,
  output     [7:0]    io_outputs_2_payload_0_0_0_6,
  output     [7:0]    io_outputs_2_payload_0_0_0_7,
  output     [7:0]    io_outputs_2_payload_0_0_0_8,
  output     [7:0]    io_outputs_2_payload_0_0_0_9,
  output     [7:0]    io_outputs_2_payload_0_0_0_10,
  output     [7:0]    io_outputs_2_payload_0_0_0_11,
  output     [7:0]    io_outputs_2_payload_0_0_0_12,
  output     [7:0]    io_outputs_2_payload_0_0_0_13,
  output     [7:0]    io_outputs_2_payload_0_0_0_14,
  output     [7:0]    io_outputs_2_payload_0_0_0_15,
  output     [7:0]    io_outputs_2_payload_0_0_1_0,
  output     [7:0]    io_outputs_2_payload_0_0_1_1,
  output     [7:0]    io_outputs_2_payload_0_0_1_2,
  output     [7:0]    io_outputs_2_payload_0_0_1_3,
  output     [7:0]    io_outputs_2_payload_0_0_1_4,
  output     [7:0]    io_outputs_2_payload_0_0_1_5,
  output     [7:0]    io_outputs_2_payload_0_0_1_6,
  output     [7:0]    io_outputs_2_payload_0_0_1_7,
  output     [7:0]    io_outputs_2_payload_0_0_1_8,
  output     [7:0]    io_outputs_2_payload_0_0_1_9,
  output     [7:0]    io_outputs_2_payload_0_0_1_10,
  output     [7:0]    io_outputs_2_payload_0_0_1_11,
  output     [7:0]    io_outputs_2_payload_0_0_1_12,
  output     [7:0]    io_outputs_2_payload_0_0_1_13,
  output     [7:0]    io_outputs_2_payload_0_0_1_14,
  output     [7:0]    io_outputs_2_payload_0_0_1_15,
  output     [7:0]    io_outputs_2_payload_0_0_2_0,
  output     [7:0]    io_outputs_2_payload_0_0_2_1,
  output     [7:0]    io_outputs_2_payload_0_0_2_2,
  output     [7:0]    io_outputs_2_payload_0_0_2_3,
  output     [7:0]    io_outputs_2_payload_0_0_2_4,
  output     [7:0]    io_outputs_2_payload_0_0_2_5,
  output     [7:0]    io_outputs_2_payload_0_0_2_6,
  output     [7:0]    io_outputs_2_payload_0_0_2_7,
  output     [7:0]    io_outputs_2_payload_0_0_2_8,
  output     [7:0]    io_outputs_2_payload_0_0_2_9,
  output     [7:0]    io_outputs_2_payload_0_0_2_10,
  output     [7:0]    io_outputs_2_payload_0_0_2_11,
  output     [7:0]    io_outputs_2_payload_0_0_2_12,
  output     [7:0]    io_outputs_2_payload_0_0_2_13,
  output     [7:0]    io_outputs_2_payload_0_0_2_14,
  output     [7:0]    io_outputs_2_payload_0_0_2_15,
  output     [7:0]    io_outputs_2_payload_0_1_0_0,
  output     [7:0]    io_outputs_2_payload_0_1_0_1,
  output     [7:0]    io_outputs_2_payload_0_1_0_2,
  output     [7:0]    io_outputs_2_payload_0_1_0_3,
  output     [7:0]    io_outputs_2_payload_0_1_0_4,
  output     [7:0]    io_outputs_2_payload_0_1_0_5,
  output     [7:0]    io_outputs_2_payload_0_1_0_6,
  output     [7:0]    io_outputs_2_payload_0_1_0_7,
  output     [7:0]    io_outputs_2_payload_0_1_0_8,
  output     [7:0]    io_outputs_2_payload_0_1_0_9,
  output     [7:0]    io_outputs_2_payload_0_1_0_10,
  output     [7:0]    io_outputs_2_payload_0_1_0_11,
  output     [7:0]    io_outputs_2_payload_0_1_0_12,
  output     [7:0]    io_outputs_2_payload_0_1_0_13,
  output     [7:0]    io_outputs_2_payload_0_1_0_14,
  output     [7:0]    io_outputs_2_payload_0_1_0_15,
  output     [7:0]    io_outputs_2_payload_0_1_1_0,
  output     [7:0]    io_outputs_2_payload_0_1_1_1,
  output     [7:0]    io_outputs_2_payload_0_1_1_2,
  output     [7:0]    io_outputs_2_payload_0_1_1_3,
  output     [7:0]    io_outputs_2_payload_0_1_1_4,
  output     [7:0]    io_outputs_2_payload_0_1_1_5,
  output     [7:0]    io_outputs_2_payload_0_1_1_6,
  output     [7:0]    io_outputs_2_payload_0_1_1_7,
  output     [7:0]    io_outputs_2_payload_0_1_1_8,
  output     [7:0]    io_outputs_2_payload_0_1_1_9,
  output     [7:0]    io_outputs_2_payload_0_1_1_10,
  output     [7:0]    io_outputs_2_payload_0_1_1_11,
  output     [7:0]    io_outputs_2_payload_0_1_1_12,
  output     [7:0]    io_outputs_2_payload_0_1_1_13,
  output     [7:0]    io_outputs_2_payload_0_1_1_14,
  output     [7:0]    io_outputs_2_payload_0_1_1_15,
  output     [7:0]    io_outputs_2_payload_0_1_2_0,
  output     [7:0]    io_outputs_2_payload_0_1_2_1,
  output     [7:0]    io_outputs_2_payload_0_1_2_2,
  output     [7:0]    io_outputs_2_payload_0_1_2_3,
  output     [7:0]    io_outputs_2_payload_0_1_2_4,
  output     [7:0]    io_outputs_2_payload_0_1_2_5,
  output     [7:0]    io_outputs_2_payload_0_1_2_6,
  output     [7:0]    io_outputs_2_payload_0_1_2_7,
  output     [7:0]    io_outputs_2_payload_0_1_2_8,
  output     [7:0]    io_outputs_2_payload_0_1_2_9,
  output     [7:0]    io_outputs_2_payload_0_1_2_10,
  output     [7:0]    io_outputs_2_payload_0_1_2_11,
  output     [7:0]    io_outputs_2_payload_0_1_2_12,
  output     [7:0]    io_outputs_2_payload_0_1_2_13,
  output     [7:0]    io_outputs_2_payload_0_1_2_14,
  output     [7:0]    io_outputs_2_payload_0_1_2_15,
  output     [7:0]    io_outputs_2_payload_0_2_0_0,
  output     [7:0]    io_outputs_2_payload_0_2_0_1,
  output     [7:0]    io_outputs_2_payload_0_2_0_2,
  output     [7:0]    io_outputs_2_payload_0_2_0_3,
  output     [7:0]    io_outputs_2_payload_0_2_0_4,
  output     [7:0]    io_outputs_2_payload_0_2_0_5,
  output     [7:0]    io_outputs_2_payload_0_2_0_6,
  output     [7:0]    io_outputs_2_payload_0_2_0_7,
  output     [7:0]    io_outputs_2_payload_0_2_0_8,
  output     [7:0]    io_outputs_2_payload_0_2_0_9,
  output     [7:0]    io_outputs_2_payload_0_2_0_10,
  output     [7:0]    io_outputs_2_payload_0_2_0_11,
  output     [7:0]    io_outputs_2_payload_0_2_0_12,
  output     [7:0]    io_outputs_2_payload_0_2_0_13,
  output     [7:0]    io_outputs_2_payload_0_2_0_14,
  output     [7:0]    io_outputs_2_payload_0_2_0_15,
  output     [7:0]    io_outputs_2_payload_0_2_1_0,
  output     [7:0]    io_outputs_2_payload_0_2_1_1,
  output     [7:0]    io_outputs_2_payload_0_2_1_2,
  output     [7:0]    io_outputs_2_payload_0_2_1_3,
  output     [7:0]    io_outputs_2_payload_0_2_1_4,
  output     [7:0]    io_outputs_2_payload_0_2_1_5,
  output     [7:0]    io_outputs_2_payload_0_2_1_6,
  output     [7:0]    io_outputs_2_payload_0_2_1_7,
  output     [7:0]    io_outputs_2_payload_0_2_1_8,
  output     [7:0]    io_outputs_2_payload_0_2_1_9,
  output     [7:0]    io_outputs_2_payload_0_2_1_10,
  output     [7:0]    io_outputs_2_payload_0_2_1_11,
  output     [7:0]    io_outputs_2_payload_0_2_1_12,
  output     [7:0]    io_outputs_2_payload_0_2_1_13,
  output     [7:0]    io_outputs_2_payload_0_2_1_14,
  output     [7:0]    io_outputs_2_payload_0_2_1_15,
  output     [7:0]    io_outputs_2_payload_0_2_2_0,
  output     [7:0]    io_outputs_2_payload_0_2_2_1,
  output     [7:0]    io_outputs_2_payload_0_2_2_2,
  output     [7:0]    io_outputs_2_payload_0_2_2_3,
  output     [7:0]    io_outputs_2_payload_0_2_2_4,
  output     [7:0]    io_outputs_2_payload_0_2_2_5,
  output     [7:0]    io_outputs_2_payload_0_2_2_6,
  output     [7:0]    io_outputs_2_payload_0_2_2_7,
  output     [7:0]    io_outputs_2_payload_0_2_2_8,
  output     [7:0]    io_outputs_2_payload_0_2_2_9,
  output     [7:0]    io_outputs_2_payload_0_2_2_10,
  output     [7:0]    io_outputs_2_payload_0_2_2_11,
  output     [7:0]    io_outputs_2_payload_0_2_2_12,
  output     [7:0]    io_outputs_2_payload_0_2_2_13,
  output     [7:0]    io_outputs_2_payload_0_2_2_14,
  output     [7:0]    io_outputs_2_payload_0_2_2_15,
  output     [7:0]    io_outputs_2_payload_1_0_0_0,
  output     [7:0]    io_outputs_2_payload_1_0_0_1,
  output     [7:0]    io_outputs_2_payload_1_0_0_2,
  output     [7:0]    io_outputs_2_payload_1_0_0_3,
  output     [7:0]    io_outputs_2_payload_1_0_0_4,
  output     [7:0]    io_outputs_2_payload_1_0_0_5,
  output     [7:0]    io_outputs_2_payload_1_0_0_6,
  output     [7:0]    io_outputs_2_payload_1_0_0_7,
  output     [7:0]    io_outputs_2_payload_1_0_0_8,
  output     [7:0]    io_outputs_2_payload_1_0_0_9,
  output     [7:0]    io_outputs_2_payload_1_0_0_10,
  output     [7:0]    io_outputs_2_payload_1_0_0_11,
  output     [7:0]    io_outputs_2_payload_1_0_0_12,
  output     [7:0]    io_outputs_2_payload_1_0_0_13,
  output     [7:0]    io_outputs_2_payload_1_0_0_14,
  output     [7:0]    io_outputs_2_payload_1_0_0_15,
  output     [7:0]    io_outputs_2_payload_1_0_1_0,
  output     [7:0]    io_outputs_2_payload_1_0_1_1,
  output     [7:0]    io_outputs_2_payload_1_0_1_2,
  output     [7:0]    io_outputs_2_payload_1_0_1_3,
  output     [7:0]    io_outputs_2_payload_1_0_1_4,
  output     [7:0]    io_outputs_2_payload_1_0_1_5,
  output     [7:0]    io_outputs_2_payload_1_0_1_6,
  output     [7:0]    io_outputs_2_payload_1_0_1_7,
  output     [7:0]    io_outputs_2_payload_1_0_1_8,
  output     [7:0]    io_outputs_2_payload_1_0_1_9,
  output     [7:0]    io_outputs_2_payload_1_0_1_10,
  output     [7:0]    io_outputs_2_payload_1_0_1_11,
  output     [7:0]    io_outputs_2_payload_1_0_1_12,
  output     [7:0]    io_outputs_2_payload_1_0_1_13,
  output     [7:0]    io_outputs_2_payload_1_0_1_14,
  output     [7:0]    io_outputs_2_payload_1_0_1_15,
  output     [7:0]    io_outputs_2_payload_1_0_2_0,
  output     [7:0]    io_outputs_2_payload_1_0_2_1,
  output     [7:0]    io_outputs_2_payload_1_0_2_2,
  output     [7:0]    io_outputs_2_payload_1_0_2_3,
  output     [7:0]    io_outputs_2_payload_1_0_2_4,
  output     [7:0]    io_outputs_2_payload_1_0_2_5,
  output     [7:0]    io_outputs_2_payload_1_0_2_6,
  output     [7:0]    io_outputs_2_payload_1_0_2_7,
  output     [7:0]    io_outputs_2_payload_1_0_2_8,
  output     [7:0]    io_outputs_2_payload_1_0_2_9,
  output     [7:0]    io_outputs_2_payload_1_0_2_10,
  output     [7:0]    io_outputs_2_payload_1_0_2_11,
  output     [7:0]    io_outputs_2_payload_1_0_2_12,
  output     [7:0]    io_outputs_2_payload_1_0_2_13,
  output     [7:0]    io_outputs_2_payload_1_0_2_14,
  output     [7:0]    io_outputs_2_payload_1_0_2_15,
  output     [7:0]    io_outputs_2_payload_1_1_0_0,
  output     [7:0]    io_outputs_2_payload_1_1_0_1,
  output     [7:0]    io_outputs_2_payload_1_1_0_2,
  output     [7:0]    io_outputs_2_payload_1_1_0_3,
  output     [7:0]    io_outputs_2_payload_1_1_0_4,
  output     [7:0]    io_outputs_2_payload_1_1_0_5,
  output     [7:0]    io_outputs_2_payload_1_1_0_6,
  output     [7:0]    io_outputs_2_payload_1_1_0_7,
  output     [7:0]    io_outputs_2_payload_1_1_0_8,
  output     [7:0]    io_outputs_2_payload_1_1_0_9,
  output     [7:0]    io_outputs_2_payload_1_1_0_10,
  output     [7:0]    io_outputs_2_payload_1_1_0_11,
  output     [7:0]    io_outputs_2_payload_1_1_0_12,
  output     [7:0]    io_outputs_2_payload_1_1_0_13,
  output     [7:0]    io_outputs_2_payload_1_1_0_14,
  output     [7:0]    io_outputs_2_payload_1_1_0_15,
  output     [7:0]    io_outputs_2_payload_1_1_1_0,
  output     [7:0]    io_outputs_2_payload_1_1_1_1,
  output     [7:0]    io_outputs_2_payload_1_1_1_2,
  output     [7:0]    io_outputs_2_payload_1_1_1_3,
  output     [7:0]    io_outputs_2_payload_1_1_1_4,
  output     [7:0]    io_outputs_2_payload_1_1_1_5,
  output     [7:0]    io_outputs_2_payload_1_1_1_6,
  output     [7:0]    io_outputs_2_payload_1_1_1_7,
  output     [7:0]    io_outputs_2_payload_1_1_1_8,
  output     [7:0]    io_outputs_2_payload_1_1_1_9,
  output     [7:0]    io_outputs_2_payload_1_1_1_10,
  output     [7:0]    io_outputs_2_payload_1_1_1_11,
  output     [7:0]    io_outputs_2_payload_1_1_1_12,
  output     [7:0]    io_outputs_2_payload_1_1_1_13,
  output     [7:0]    io_outputs_2_payload_1_1_1_14,
  output     [7:0]    io_outputs_2_payload_1_1_1_15,
  output     [7:0]    io_outputs_2_payload_1_1_2_0,
  output     [7:0]    io_outputs_2_payload_1_1_2_1,
  output     [7:0]    io_outputs_2_payload_1_1_2_2,
  output     [7:0]    io_outputs_2_payload_1_1_2_3,
  output     [7:0]    io_outputs_2_payload_1_1_2_4,
  output     [7:0]    io_outputs_2_payload_1_1_2_5,
  output     [7:0]    io_outputs_2_payload_1_1_2_6,
  output     [7:0]    io_outputs_2_payload_1_1_2_7,
  output     [7:0]    io_outputs_2_payload_1_1_2_8,
  output     [7:0]    io_outputs_2_payload_1_1_2_9,
  output     [7:0]    io_outputs_2_payload_1_1_2_10,
  output     [7:0]    io_outputs_2_payload_1_1_2_11,
  output     [7:0]    io_outputs_2_payload_1_1_2_12,
  output     [7:0]    io_outputs_2_payload_1_1_2_13,
  output     [7:0]    io_outputs_2_payload_1_1_2_14,
  output     [7:0]    io_outputs_2_payload_1_1_2_15,
  output     [7:0]    io_outputs_2_payload_1_2_0_0,
  output     [7:0]    io_outputs_2_payload_1_2_0_1,
  output     [7:0]    io_outputs_2_payload_1_2_0_2,
  output     [7:0]    io_outputs_2_payload_1_2_0_3,
  output     [7:0]    io_outputs_2_payload_1_2_0_4,
  output     [7:0]    io_outputs_2_payload_1_2_0_5,
  output     [7:0]    io_outputs_2_payload_1_2_0_6,
  output     [7:0]    io_outputs_2_payload_1_2_0_7,
  output     [7:0]    io_outputs_2_payload_1_2_0_8,
  output     [7:0]    io_outputs_2_payload_1_2_0_9,
  output     [7:0]    io_outputs_2_payload_1_2_0_10,
  output     [7:0]    io_outputs_2_payload_1_2_0_11,
  output     [7:0]    io_outputs_2_payload_1_2_0_12,
  output     [7:0]    io_outputs_2_payload_1_2_0_13,
  output     [7:0]    io_outputs_2_payload_1_2_0_14,
  output     [7:0]    io_outputs_2_payload_1_2_0_15,
  output     [7:0]    io_outputs_2_payload_1_2_1_0,
  output     [7:0]    io_outputs_2_payload_1_2_1_1,
  output     [7:0]    io_outputs_2_payload_1_2_1_2,
  output     [7:0]    io_outputs_2_payload_1_2_1_3,
  output     [7:0]    io_outputs_2_payload_1_2_1_4,
  output     [7:0]    io_outputs_2_payload_1_2_1_5,
  output     [7:0]    io_outputs_2_payload_1_2_1_6,
  output     [7:0]    io_outputs_2_payload_1_2_1_7,
  output     [7:0]    io_outputs_2_payload_1_2_1_8,
  output     [7:0]    io_outputs_2_payload_1_2_1_9,
  output     [7:0]    io_outputs_2_payload_1_2_1_10,
  output     [7:0]    io_outputs_2_payload_1_2_1_11,
  output     [7:0]    io_outputs_2_payload_1_2_1_12,
  output     [7:0]    io_outputs_2_payload_1_2_1_13,
  output     [7:0]    io_outputs_2_payload_1_2_1_14,
  output     [7:0]    io_outputs_2_payload_1_2_1_15,
  output     [7:0]    io_outputs_2_payload_1_2_2_0,
  output     [7:0]    io_outputs_2_payload_1_2_2_1,
  output     [7:0]    io_outputs_2_payload_1_2_2_2,
  output     [7:0]    io_outputs_2_payload_1_2_2_3,
  output     [7:0]    io_outputs_2_payload_1_2_2_4,
  output     [7:0]    io_outputs_2_payload_1_2_2_5,
  output     [7:0]    io_outputs_2_payload_1_2_2_6,
  output     [7:0]    io_outputs_2_payload_1_2_2_7,
  output     [7:0]    io_outputs_2_payload_1_2_2_8,
  output     [7:0]    io_outputs_2_payload_1_2_2_9,
  output     [7:0]    io_outputs_2_payload_1_2_2_10,
  output     [7:0]    io_outputs_2_payload_1_2_2_11,
  output     [7:0]    io_outputs_2_payload_1_2_2_12,
  output     [7:0]    io_outputs_2_payload_1_2_2_13,
  output     [7:0]    io_outputs_2_payload_1_2_2_14,
  output     [7:0]    io_outputs_2_payload_1_2_2_15,
  output reg          io_outputs_3_valid,
  input               io_outputs_3_ready,
  output     [7:0]    io_outputs_3_payload_0_0_0_0,
  output     [7:0]    io_outputs_3_payload_0_0_0_1,
  output     [7:0]    io_outputs_3_payload_0_0_0_2,
  output     [7:0]    io_outputs_3_payload_0_0_0_3,
  output     [7:0]    io_outputs_3_payload_0_0_0_4,
  output     [7:0]    io_outputs_3_payload_0_0_0_5,
  output     [7:0]    io_outputs_3_payload_0_0_0_6,
  output     [7:0]    io_outputs_3_payload_0_0_0_7,
  output     [7:0]    io_outputs_3_payload_0_0_0_8,
  output     [7:0]    io_outputs_3_payload_0_0_0_9,
  output     [7:0]    io_outputs_3_payload_0_0_0_10,
  output     [7:0]    io_outputs_3_payload_0_0_0_11,
  output     [7:0]    io_outputs_3_payload_0_0_0_12,
  output     [7:0]    io_outputs_3_payload_0_0_0_13,
  output     [7:0]    io_outputs_3_payload_0_0_0_14,
  output     [7:0]    io_outputs_3_payload_0_0_0_15,
  output     [7:0]    io_outputs_3_payload_0_0_1_0,
  output     [7:0]    io_outputs_3_payload_0_0_1_1,
  output     [7:0]    io_outputs_3_payload_0_0_1_2,
  output     [7:0]    io_outputs_3_payload_0_0_1_3,
  output     [7:0]    io_outputs_3_payload_0_0_1_4,
  output     [7:0]    io_outputs_3_payload_0_0_1_5,
  output     [7:0]    io_outputs_3_payload_0_0_1_6,
  output     [7:0]    io_outputs_3_payload_0_0_1_7,
  output     [7:0]    io_outputs_3_payload_0_0_1_8,
  output     [7:0]    io_outputs_3_payload_0_0_1_9,
  output     [7:0]    io_outputs_3_payload_0_0_1_10,
  output     [7:0]    io_outputs_3_payload_0_0_1_11,
  output     [7:0]    io_outputs_3_payload_0_0_1_12,
  output     [7:0]    io_outputs_3_payload_0_0_1_13,
  output     [7:0]    io_outputs_3_payload_0_0_1_14,
  output     [7:0]    io_outputs_3_payload_0_0_1_15,
  output     [7:0]    io_outputs_3_payload_0_0_2_0,
  output     [7:0]    io_outputs_3_payload_0_0_2_1,
  output     [7:0]    io_outputs_3_payload_0_0_2_2,
  output     [7:0]    io_outputs_3_payload_0_0_2_3,
  output     [7:0]    io_outputs_3_payload_0_0_2_4,
  output     [7:0]    io_outputs_3_payload_0_0_2_5,
  output     [7:0]    io_outputs_3_payload_0_0_2_6,
  output     [7:0]    io_outputs_3_payload_0_0_2_7,
  output     [7:0]    io_outputs_3_payload_0_0_2_8,
  output     [7:0]    io_outputs_3_payload_0_0_2_9,
  output     [7:0]    io_outputs_3_payload_0_0_2_10,
  output     [7:0]    io_outputs_3_payload_0_0_2_11,
  output     [7:0]    io_outputs_3_payload_0_0_2_12,
  output     [7:0]    io_outputs_3_payload_0_0_2_13,
  output     [7:0]    io_outputs_3_payload_0_0_2_14,
  output     [7:0]    io_outputs_3_payload_0_0_2_15,
  output     [7:0]    io_outputs_3_payload_0_1_0_0,
  output     [7:0]    io_outputs_3_payload_0_1_0_1,
  output     [7:0]    io_outputs_3_payload_0_1_0_2,
  output     [7:0]    io_outputs_3_payload_0_1_0_3,
  output     [7:0]    io_outputs_3_payload_0_1_0_4,
  output     [7:0]    io_outputs_3_payload_0_1_0_5,
  output     [7:0]    io_outputs_3_payload_0_1_0_6,
  output     [7:0]    io_outputs_3_payload_0_1_0_7,
  output     [7:0]    io_outputs_3_payload_0_1_0_8,
  output     [7:0]    io_outputs_3_payload_0_1_0_9,
  output     [7:0]    io_outputs_3_payload_0_1_0_10,
  output     [7:0]    io_outputs_3_payload_0_1_0_11,
  output     [7:0]    io_outputs_3_payload_0_1_0_12,
  output     [7:0]    io_outputs_3_payload_0_1_0_13,
  output     [7:0]    io_outputs_3_payload_0_1_0_14,
  output     [7:0]    io_outputs_3_payload_0_1_0_15,
  output     [7:0]    io_outputs_3_payload_0_1_1_0,
  output     [7:0]    io_outputs_3_payload_0_1_1_1,
  output     [7:0]    io_outputs_3_payload_0_1_1_2,
  output     [7:0]    io_outputs_3_payload_0_1_1_3,
  output     [7:0]    io_outputs_3_payload_0_1_1_4,
  output     [7:0]    io_outputs_3_payload_0_1_1_5,
  output     [7:0]    io_outputs_3_payload_0_1_1_6,
  output     [7:0]    io_outputs_3_payload_0_1_1_7,
  output     [7:0]    io_outputs_3_payload_0_1_1_8,
  output     [7:0]    io_outputs_3_payload_0_1_1_9,
  output     [7:0]    io_outputs_3_payload_0_1_1_10,
  output     [7:0]    io_outputs_3_payload_0_1_1_11,
  output     [7:0]    io_outputs_3_payload_0_1_1_12,
  output     [7:0]    io_outputs_3_payload_0_1_1_13,
  output     [7:0]    io_outputs_3_payload_0_1_1_14,
  output     [7:0]    io_outputs_3_payload_0_1_1_15,
  output     [7:0]    io_outputs_3_payload_0_1_2_0,
  output     [7:0]    io_outputs_3_payload_0_1_2_1,
  output     [7:0]    io_outputs_3_payload_0_1_2_2,
  output     [7:0]    io_outputs_3_payload_0_1_2_3,
  output     [7:0]    io_outputs_3_payload_0_1_2_4,
  output     [7:0]    io_outputs_3_payload_0_1_2_5,
  output     [7:0]    io_outputs_3_payload_0_1_2_6,
  output     [7:0]    io_outputs_3_payload_0_1_2_7,
  output     [7:0]    io_outputs_3_payload_0_1_2_8,
  output     [7:0]    io_outputs_3_payload_0_1_2_9,
  output     [7:0]    io_outputs_3_payload_0_1_2_10,
  output     [7:0]    io_outputs_3_payload_0_1_2_11,
  output     [7:0]    io_outputs_3_payload_0_1_2_12,
  output     [7:0]    io_outputs_3_payload_0_1_2_13,
  output     [7:0]    io_outputs_3_payload_0_1_2_14,
  output     [7:0]    io_outputs_3_payload_0_1_2_15,
  output     [7:0]    io_outputs_3_payload_0_2_0_0,
  output     [7:0]    io_outputs_3_payload_0_2_0_1,
  output     [7:0]    io_outputs_3_payload_0_2_0_2,
  output     [7:0]    io_outputs_3_payload_0_2_0_3,
  output     [7:0]    io_outputs_3_payload_0_2_0_4,
  output     [7:0]    io_outputs_3_payload_0_2_0_5,
  output     [7:0]    io_outputs_3_payload_0_2_0_6,
  output     [7:0]    io_outputs_3_payload_0_2_0_7,
  output     [7:0]    io_outputs_3_payload_0_2_0_8,
  output     [7:0]    io_outputs_3_payload_0_2_0_9,
  output     [7:0]    io_outputs_3_payload_0_2_0_10,
  output     [7:0]    io_outputs_3_payload_0_2_0_11,
  output     [7:0]    io_outputs_3_payload_0_2_0_12,
  output     [7:0]    io_outputs_3_payload_0_2_0_13,
  output     [7:0]    io_outputs_3_payload_0_2_0_14,
  output     [7:0]    io_outputs_3_payload_0_2_0_15,
  output     [7:0]    io_outputs_3_payload_0_2_1_0,
  output     [7:0]    io_outputs_3_payload_0_2_1_1,
  output     [7:0]    io_outputs_3_payload_0_2_1_2,
  output     [7:0]    io_outputs_3_payload_0_2_1_3,
  output     [7:0]    io_outputs_3_payload_0_2_1_4,
  output     [7:0]    io_outputs_3_payload_0_2_1_5,
  output     [7:0]    io_outputs_3_payload_0_2_1_6,
  output     [7:0]    io_outputs_3_payload_0_2_1_7,
  output     [7:0]    io_outputs_3_payload_0_2_1_8,
  output     [7:0]    io_outputs_3_payload_0_2_1_9,
  output     [7:0]    io_outputs_3_payload_0_2_1_10,
  output     [7:0]    io_outputs_3_payload_0_2_1_11,
  output     [7:0]    io_outputs_3_payload_0_2_1_12,
  output     [7:0]    io_outputs_3_payload_0_2_1_13,
  output     [7:0]    io_outputs_3_payload_0_2_1_14,
  output     [7:0]    io_outputs_3_payload_0_2_1_15,
  output     [7:0]    io_outputs_3_payload_0_2_2_0,
  output     [7:0]    io_outputs_3_payload_0_2_2_1,
  output     [7:0]    io_outputs_3_payload_0_2_2_2,
  output     [7:0]    io_outputs_3_payload_0_2_2_3,
  output     [7:0]    io_outputs_3_payload_0_2_2_4,
  output     [7:0]    io_outputs_3_payload_0_2_2_5,
  output     [7:0]    io_outputs_3_payload_0_2_2_6,
  output     [7:0]    io_outputs_3_payload_0_2_2_7,
  output     [7:0]    io_outputs_3_payload_0_2_2_8,
  output     [7:0]    io_outputs_3_payload_0_2_2_9,
  output     [7:0]    io_outputs_3_payload_0_2_2_10,
  output     [7:0]    io_outputs_3_payload_0_2_2_11,
  output     [7:0]    io_outputs_3_payload_0_2_2_12,
  output     [7:0]    io_outputs_3_payload_0_2_2_13,
  output     [7:0]    io_outputs_3_payload_0_2_2_14,
  output     [7:0]    io_outputs_3_payload_0_2_2_15,
  output     [7:0]    io_outputs_3_payload_1_0_0_0,
  output     [7:0]    io_outputs_3_payload_1_0_0_1,
  output     [7:0]    io_outputs_3_payload_1_0_0_2,
  output     [7:0]    io_outputs_3_payload_1_0_0_3,
  output     [7:0]    io_outputs_3_payload_1_0_0_4,
  output     [7:0]    io_outputs_3_payload_1_0_0_5,
  output     [7:0]    io_outputs_3_payload_1_0_0_6,
  output     [7:0]    io_outputs_3_payload_1_0_0_7,
  output     [7:0]    io_outputs_3_payload_1_0_0_8,
  output     [7:0]    io_outputs_3_payload_1_0_0_9,
  output     [7:0]    io_outputs_3_payload_1_0_0_10,
  output     [7:0]    io_outputs_3_payload_1_0_0_11,
  output     [7:0]    io_outputs_3_payload_1_0_0_12,
  output     [7:0]    io_outputs_3_payload_1_0_0_13,
  output     [7:0]    io_outputs_3_payload_1_0_0_14,
  output     [7:0]    io_outputs_3_payload_1_0_0_15,
  output     [7:0]    io_outputs_3_payload_1_0_1_0,
  output     [7:0]    io_outputs_3_payload_1_0_1_1,
  output     [7:0]    io_outputs_3_payload_1_0_1_2,
  output     [7:0]    io_outputs_3_payload_1_0_1_3,
  output     [7:0]    io_outputs_3_payload_1_0_1_4,
  output     [7:0]    io_outputs_3_payload_1_0_1_5,
  output     [7:0]    io_outputs_3_payload_1_0_1_6,
  output     [7:0]    io_outputs_3_payload_1_0_1_7,
  output     [7:0]    io_outputs_3_payload_1_0_1_8,
  output     [7:0]    io_outputs_3_payload_1_0_1_9,
  output     [7:0]    io_outputs_3_payload_1_0_1_10,
  output     [7:0]    io_outputs_3_payload_1_0_1_11,
  output     [7:0]    io_outputs_3_payload_1_0_1_12,
  output     [7:0]    io_outputs_3_payload_1_0_1_13,
  output     [7:0]    io_outputs_3_payload_1_0_1_14,
  output     [7:0]    io_outputs_3_payload_1_0_1_15,
  output     [7:0]    io_outputs_3_payload_1_0_2_0,
  output     [7:0]    io_outputs_3_payload_1_0_2_1,
  output     [7:0]    io_outputs_3_payload_1_0_2_2,
  output     [7:0]    io_outputs_3_payload_1_0_2_3,
  output     [7:0]    io_outputs_3_payload_1_0_2_4,
  output     [7:0]    io_outputs_3_payload_1_0_2_5,
  output     [7:0]    io_outputs_3_payload_1_0_2_6,
  output     [7:0]    io_outputs_3_payload_1_0_2_7,
  output     [7:0]    io_outputs_3_payload_1_0_2_8,
  output     [7:0]    io_outputs_3_payload_1_0_2_9,
  output     [7:0]    io_outputs_3_payload_1_0_2_10,
  output     [7:0]    io_outputs_3_payload_1_0_2_11,
  output     [7:0]    io_outputs_3_payload_1_0_2_12,
  output     [7:0]    io_outputs_3_payload_1_0_2_13,
  output     [7:0]    io_outputs_3_payload_1_0_2_14,
  output     [7:0]    io_outputs_3_payload_1_0_2_15,
  output     [7:0]    io_outputs_3_payload_1_1_0_0,
  output     [7:0]    io_outputs_3_payload_1_1_0_1,
  output     [7:0]    io_outputs_3_payload_1_1_0_2,
  output     [7:0]    io_outputs_3_payload_1_1_0_3,
  output     [7:0]    io_outputs_3_payload_1_1_0_4,
  output     [7:0]    io_outputs_3_payload_1_1_0_5,
  output     [7:0]    io_outputs_3_payload_1_1_0_6,
  output     [7:0]    io_outputs_3_payload_1_1_0_7,
  output     [7:0]    io_outputs_3_payload_1_1_0_8,
  output     [7:0]    io_outputs_3_payload_1_1_0_9,
  output     [7:0]    io_outputs_3_payload_1_1_0_10,
  output     [7:0]    io_outputs_3_payload_1_1_0_11,
  output     [7:0]    io_outputs_3_payload_1_1_0_12,
  output     [7:0]    io_outputs_3_payload_1_1_0_13,
  output     [7:0]    io_outputs_3_payload_1_1_0_14,
  output     [7:0]    io_outputs_3_payload_1_1_0_15,
  output     [7:0]    io_outputs_3_payload_1_1_1_0,
  output     [7:0]    io_outputs_3_payload_1_1_1_1,
  output     [7:0]    io_outputs_3_payload_1_1_1_2,
  output     [7:0]    io_outputs_3_payload_1_1_1_3,
  output     [7:0]    io_outputs_3_payload_1_1_1_4,
  output     [7:0]    io_outputs_3_payload_1_1_1_5,
  output     [7:0]    io_outputs_3_payload_1_1_1_6,
  output     [7:0]    io_outputs_3_payload_1_1_1_7,
  output     [7:0]    io_outputs_3_payload_1_1_1_8,
  output     [7:0]    io_outputs_3_payload_1_1_1_9,
  output     [7:0]    io_outputs_3_payload_1_1_1_10,
  output     [7:0]    io_outputs_3_payload_1_1_1_11,
  output     [7:0]    io_outputs_3_payload_1_1_1_12,
  output     [7:0]    io_outputs_3_payload_1_1_1_13,
  output     [7:0]    io_outputs_3_payload_1_1_1_14,
  output     [7:0]    io_outputs_3_payload_1_1_1_15,
  output     [7:0]    io_outputs_3_payload_1_1_2_0,
  output     [7:0]    io_outputs_3_payload_1_1_2_1,
  output     [7:0]    io_outputs_3_payload_1_1_2_2,
  output     [7:0]    io_outputs_3_payload_1_1_2_3,
  output     [7:0]    io_outputs_3_payload_1_1_2_4,
  output     [7:0]    io_outputs_3_payload_1_1_2_5,
  output     [7:0]    io_outputs_3_payload_1_1_2_6,
  output     [7:0]    io_outputs_3_payload_1_1_2_7,
  output     [7:0]    io_outputs_3_payload_1_1_2_8,
  output     [7:0]    io_outputs_3_payload_1_1_2_9,
  output     [7:0]    io_outputs_3_payload_1_1_2_10,
  output     [7:0]    io_outputs_3_payload_1_1_2_11,
  output     [7:0]    io_outputs_3_payload_1_1_2_12,
  output     [7:0]    io_outputs_3_payload_1_1_2_13,
  output     [7:0]    io_outputs_3_payload_1_1_2_14,
  output     [7:0]    io_outputs_3_payload_1_1_2_15,
  output     [7:0]    io_outputs_3_payload_1_2_0_0,
  output     [7:0]    io_outputs_3_payload_1_2_0_1,
  output     [7:0]    io_outputs_3_payload_1_2_0_2,
  output     [7:0]    io_outputs_3_payload_1_2_0_3,
  output     [7:0]    io_outputs_3_payload_1_2_0_4,
  output     [7:0]    io_outputs_3_payload_1_2_0_5,
  output     [7:0]    io_outputs_3_payload_1_2_0_6,
  output     [7:0]    io_outputs_3_payload_1_2_0_7,
  output     [7:0]    io_outputs_3_payload_1_2_0_8,
  output     [7:0]    io_outputs_3_payload_1_2_0_9,
  output     [7:0]    io_outputs_3_payload_1_2_0_10,
  output     [7:0]    io_outputs_3_payload_1_2_0_11,
  output     [7:0]    io_outputs_3_payload_1_2_0_12,
  output     [7:0]    io_outputs_3_payload_1_2_0_13,
  output     [7:0]    io_outputs_3_payload_1_2_0_14,
  output     [7:0]    io_outputs_3_payload_1_2_0_15,
  output     [7:0]    io_outputs_3_payload_1_2_1_0,
  output     [7:0]    io_outputs_3_payload_1_2_1_1,
  output     [7:0]    io_outputs_3_payload_1_2_1_2,
  output     [7:0]    io_outputs_3_payload_1_2_1_3,
  output     [7:0]    io_outputs_3_payload_1_2_1_4,
  output     [7:0]    io_outputs_3_payload_1_2_1_5,
  output     [7:0]    io_outputs_3_payload_1_2_1_6,
  output     [7:0]    io_outputs_3_payload_1_2_1_7,
  output     [7:0]    io_outputs_3_payload_1_2_1_8,
  output     [7:0]    io_outputs_3_payload_1_2_1_9,
  output     [7:0]    io_outputs_3_payload_1_2_1_10,
  output     [7:0]    io_outputs_3_payload_1_2_1_11,
  output     [7:0]    io_outputs_3_payload_1_2_1_12,
  output     [7:0]    io_outputs_3_payload_1_2_1_13,
  output     [7:0]    io_outputs_3_payload_1_2_1_14,
  output     [7:0]    io_outputs_3_payload_1_2_1_15,
  output     [7:0]    io_outputs_3_payload_1_2_2_0,
  output     [7:0]    io_outputs_3_payload_1_2_2_1,
  output     [7:0]    io_outputs_3_payload_1_2_2_2,
  output     [7:0]    io_outputs_3_payload_1_2_2_3,
  output     [7:0]    io_outputs_3_payload_1_2_2_4,
  output     [7:0]    io_outputs_3_payload_1_2_2_5,
  output     [7:0]    io_outputs_3_payload_1_2_2_6,
  output     [7:0]    io_outputs_3_payload_1_2_2_7,
  output     [7:0]    io_outputs_3_payload_1_2_2_8,
  output     [7:0]    io_outputs_3_payload_1_2_2_9,
  output     [7:0]    io_outputs_3_payload_1_2_2_10,
  output     [7:0]    io_outputs_3_payload_1_2_2_11,
  output     [7:0]    io_outputs_3_payload_1_2_2_12,
  output     [7:0]    io_outputs_3_payload_1_2_2_13,
  output     [7:0]    io_outputs_3_payload_1_2_2_14,
  output     [7:0]    io_outputs_3_payload_1_2_2_15,
  output reg          io_outputs_4_valid,
  input               io_outputs_4_ready,
  output     [7:0]    io_outputs_4_payload_0_0_0_0,
  output     [7:0]    io_outputs_4_payload_0_0_0_1,
  output     [7:0]    io_outputs_4_payload_0_0_0_2,
  output     [7:0]    io_outputs_4_payload_0_0_0_3,
  output     [7:0]    io_outputs_4_payload_0_0_0_4,
  output     [7:0]    io_outputs_4_payload_0_0_0_5,
  output     [7:0]    io_outputs_4_payload_0_0_0_6,
  output     [7:0]    io_outputs_4_payload_0_0_0_7,
  output     [7:0]    io_outputs_4_payload_0_0_0_8,
  output     [7:0]    io_outputs_4_payload_0_0_0_9,
  output     [7:0]    io_outputs_4_payload_0_0_0_10,
  output     [7:0]    io_outputs_4_payload_0_0_0_11,
  output     [7:0]    io_outputs_4_payload_0_0_0_12,
  output     [7:0]    io_outputs_4_payload_0_0_0_13,
  output     [7:0]    io_outputs_4_payload_0_0_0_14,
  output     [7:0]    io_outputs_4_payload_0_0_0_15,
  output     [7:0]    io_outputs_4_payload_0_0_1_0,
  output     [7:0]    io_outputs_4_payload_0_0_1_1,
  output     [7:0]    io_outputs_4_payload_0_0_1_2,
  output     [7:0]    io_outputs_4_payload_0_0_1_3,
  output     [7:0]    io_outputs_4_payload_0_0_1_4,
  output     [7:0]    io_outputs_4_payload_0_0_1_5,
  output     [7:0]    io_outputs_4_payload_0_0_1_6,
  output     [7:0]    io_outputs_4_payload_0_0_1_7,
  output     [7:0]    io_outputs_4_payload_0_0_1_8,
  output     [7:0]    io_outputs_4_payload_0_0_1_9,
  output     [7:0]    io_outputs_4_payload_0_0_1_10,
  output     [7:0]    io_outputs_4_payload_0_0_1_11,
  output     [7:0]    io_outputs_4_payload_0_0_1_12,
  output     [7:0]    io_outputs_4_payload_0_0_1_13,
  output     [7:0]    io_outputs_4_payload_0_0_1_14,
  output     [7:0]    io_outputs_4_payload_0_0_1_15,
  output     [7:0]    io_outputs_4_payload_0_0_2_0,
  output     [7:0]    io_outputs_4_payload_0_0_2_1,
  output     [7:0]    io_outputs_4_payload_0_0_2_2,
  output     [7:0]    io_outputs_4_payload_0_0_2_3,
  output     [7:0]    io_outputs_4_payload_0_0_2_4,
  output     [7:0]    io_outputs_4_payload_0_0_2_5,
  output     [7:0]    io_outputs_4_payload_0_0_2_6,
  output     [7:0]    io_outputs_4_payload_0_0_2_7,
  output     [7:0]    io_outputs_4_payload_0_0_2_8,
  output     [7:0]    io_outputs_4_payload_0_0_2_9,
  output     [7:0]    io_outputs_4_payload_0_0_2_10,
  output     [7:0]    io_outputs_4_payload_0_0_2_11,
  output     [7:0]    io_outputs_4_payload_0_0_2_12,
  output     [7:0]    io_outputs_4_payload_0_0_2_13,
  output     [7:0]    io_outputs_4_payload_0_0_2_14,
  output     [7:0]    io_outputs_4_payload_0_0_2_15,
  output     [7:0]    io_outputs_4_payload_0_1_0_0,
  output     [7:0]    io_outputs_4_payload_0_1_0_1,
  output     [7:0]    io_outputs_4_payload_0_1_0_2,
  output     [7:0]    io_outputs_4_payload_0_1_0_3,
  output     [7:0]    io_outputs_4_payload_0_1_0_4,
  output     [7:0]    io_outputs_4_payload_0_1_0_5,
  output     [7:0]    io_outputs_4_payload_0_1_0_6,
  output     [7:0]    io_outputs_4_payload_0_1_0_7,
  output     [7:0]    io_outputs_4_payload_0_1_0_8,
  output     [7:0]    io_outputs_4_payload_0_1_0_9,
  output     [7:0]    io_outputs_4_payload_0_1_0_10,
  output     [7:0]    io_outputs_4_payload_0_1_0_11,
  output     [7:0]    io_outputs_4_payload_0_1_0_12,
  output     [7:0]    io_outputs_4_payload_0_1_0_13,
  output     [7:0]    io_outputs_4_payload_0_1_0_14,
  output     [7:0]    io_outputs_4_payload_0_1_0_15,
  output     [7:0]    io_outputs_4_payload_0_1_1_0,
  output     [7:0]    io_outputs_4_payload_0_1_1_1,
  output     [7:0]    io_outputs_4_payload_0_1_1_2,
  output     [7:0]    io_outputs_4_payload_0_1_1_3,
  output     [7:0]    io_outputs_4_payload_0_1_1_4,
  output     [7:0]    io_outputs_4_payload_0_1_1_5,
  output     [7:0]    io_outputs_4_payload_0_1_1_6,
  output     [7:0]    io_outputs_4_payload_0_1_1_7,
  output     [7:0]    io_outputs_4_payload_0_1_1_8,
  output     [7:0]    io_outputs_4_payload_0_1_1_9,
  output     [7:0]    io_outputs_4_payload_0_1_1_10,
  output     [7:0]    io_outputs_4_payload_0_1_1_11,
  output     [7:0]    io_outputs_4_payload_0_1_1_12,
  output     [7:0]    io_outputs_4_payload_0_1_1_13,
  output     [7:0]    io_outputs_4_payload_0_1_1_14,
  output     [7:0]    io_outputs_4_payload_0_1_1_15,
  output     [7:0]    io_outputs_4_payload_0_1_2_0,
  output     [7:0]    io_outputs_4_payload_0_1_2_1,
  output     [7:0]    io_outputs_4_payload_0_1_2_2,
  output     [7:0]    io_outputs_4_payload_0_1_2_3,
  output     [7:0]    io_outputs_4_payload_0_1_2_4,
  output     [7:0]    io_outputs_4_payload_0_1_2_5,
  output     [7:0]    io_outputs_4_payload_0_1_2_6,
  output     [7:0]    io_outputs_4_payload_0_1_2_7,
  output     [7:0]    io_outputs_4_payload_0_1_2_8,
  output     [7:0]    io_outputs_4_payload_0_1_2_9,
  output     [7:0]    io_outputs_4_payload_0_1_2_10,
  output     [7:0]    io_outputs_4_payload_0_1_2_11,
  output     [7:0]    io_outputs_4_payload_0_1_2_12,
  output     [7:0]    io_outputs_4_payload_0_1_2_13,
  output     [7:0]    io_outputs_4_payload_0_1_2_14,
  output     [7:0]    io_outputs_4_payload_0_1_2_15,
  output     [7:0]    io_outputs_4_payload_0_2_0_0,
  output     [7:0]    io_outputs_4_payload_0_2_0_1,
  output     [7:0]    io_outputs_4_payload_0_2_0_2,
  output     [7:0]    io_outputs_4_payload_0_2_0_3,
  output     [7:0]    io_outputs_4_payload_0_2_0_4,
  output     [7:0]    io_outputs_4_payload_0_2_0_5,
  output     [7:0]    io_outputs_4_payload_0_2_0_6,
  output     [7:0]    io_outputs_4_payload_0_2_0_7,
  output     [7:0]    io_outputs_4_payload_0_2_0_8,
  output     [7:0]    io_outputs_4_payload_0_2_0_9,
  output     [7:0]    io_outputs_4_payload_0_2_0_10,
  output     [7:0]    io_outputs_4_payload_0_2_0_11,
  output     [7:0]    io_outputs_4_payload_0_2_0_12,
  output     [7:0]    io_outputs_4_payload_0_2_0_13,
  output     [7:0]    io_outputs_4_payload_0_2_0_14,
  output     [7:0]    io_outputs_4_payload_0_2_0_15,
  output     [7:0]    io_outputs_4_payload_0_2_1_0,
  output     [7:0]    io_outputs_4_payload_0_2_1_1,
  output     [7:0]    io_outputs_4_payload_0_2_1_2,
  output     [7:0]    io_outputs_4_payload_0_2_1_3,
  output     [7:0]    io_outputs_4_payload_0_2_1_4,
  output     [7:0]    io_outputs_4_payload_0_2_1_5,
  output     [7:0]    io_outputs_4_payload_0_2_1_6,
  output     [7:0]    io_outputs_4_payload_0_2_1_7,
  output     [7:0]    io_outputs_4_payload_0_2_1_8,
  output     [7:0]    io_outputs_4_payload_0_2_1_9,
  output     [7:0]    io_outputs_4_payload_0_2_1_10,
  output     [7:0]    io_outputs_4_payload_0_2_1_11,
  output     [7:0]    io_outputs_4_payload_0_2_1_12,
  output     [7:0]    io_outputs_4_payload_0_2_1_13,
  output     [7:0]    io_outputs_4_payload_0_2_1_14,
  output     [7:0]    io_outputs_4_payload_0_2_1_15,
  output     [7:0]    io_outputs_4_payload_0_2_2_0,
  output     [7:0]    io_outputs_4_payload_0_2_2_1,
  output     [7:0]    io_outputs_4_payload_0_2_2_2,
  output     [7:0]    io_outputs_4_payload_0_2_2_3,
  output     [7:0]    io_outputs_4_payload_0_2_2_4,
  output     [7:0]    io_outputs_4_payload_0_2_2_5,
  output     [7:0]    io_outputs_4_payload_0_2_2_6,
  output     [7:0]    io_outputs_4_payload_0_2_2_7,
  output     [7:0]    io_outputs_4_payload_0_2_2_8,
  output     [7:0]    io_outputs_4_payload_0_2_2_9,
  output     [7:0]    io_outputs_4_payload_0_2_2_10,
  output     [7:0]    io_outputs_4_payload_0_2_2_11,
  output     [7:0]    io_outputs_4_payload_0_2_2_12,
  output     [7:0]    io_outputs_4_payload_0_2_2_13,
  output     [7:0]    io_outputs_4_payload_0_2_2_14,
  output     [7:0]    io_outputs_4_payload_0_2_2_15,
  output     [7:0]    io_outputs_4_payload_1_0_0_0,
  output     [7:0]    io_outputs_4_payload_1_0_0_1,
  output     [7:0]    io_outputs_4_payload_1_0_0_2,
  output     [7:0]    io_outputs_4_payload_1_0_0_3,
  output     [7:0]    io_outputs_4_payload_1_0_0_4,
  output     [7:0]    io_outputs_4_payload_1_0_0_5,
  output     [7:0]    io_outputs_4_payload_1_0_0_6,
  output     [7:0]    io_outputs_4_payload_1_0_0_7,
  output     [7:0]    io_outputs_4_payload_1_0_0_8,
  output     [7:0]    io_outputs_4_payload_1_0_0_9,
  output     [7:0]    io_outputs_4_payload_1_0_0_10,
  output     [7:0]    io_outputs_4_payload_1_0_0_11,
  output     [7:0]    io_outputs_4_payload_1_0_0_12,
  output     [7:0]    io_outputs_4_payload_1_0_0_13,
  output     [7:0]    io_outputs_4_payload_1_0_0_14,
  output     [7:0]    io_outputs_4_payload_1_0_0_15,
  output     [7:0]    io_outputs_4_payload_1_0_1_0,
  output     [7:0]    io_outputs_4_payload_1_0_1_1,
  output     [7:0]    io_outputs_4_payload_1_0_1_2,
  output     [7:0]    io_outputs_4_payload_1_0_1_3,
  output     [7:0]    io_outputs_4_payload_1_0_1_4,
  output     [7:0]    io_outputs_4_payload_1_0_1_5,
  output     [7:0]    io_outputs_4_payload_1_0_1_6,
  output     [7:0]    io_outputs_4_payload_1_0_1_7,
  output     [7:0]    io_outputs_4_payload_1_0_1_8,
  output     [7:0]    io_outputs_4_payload_1_0_1_9,
  output     [7:0]    io_outputs_4_payload_1_0_1_10,
  output     [7:0]    io_outputs_4_payload_1_0_1_11,
  output     [7:0]    io_outputs_4_payload_1_0_1_12,
  output     [7:0]    io_outputs_4_payload_1_0_1_13,
  output     [7:0]    io_outputs_4_payload_1_0_1_14,
  output     [7:0]    io_outputs_4_payload_1_0_1_15,
  output     [7:0]    io_outputs_4_payload_1_0_2_0,
  output     [7:0]    io_outputs_4_payload_1_0_2_1,
  output     [7:0]    io_outputs_4_payload_1_0_2_2,
  output     [7:0]    io_outputs_4_payload_1_0_2_3,
  output     [7:0]    io_outputs_4_payload_1_0_2_4,
  output     [7:0]    io_outputs_4_payload_1_0_2_5,
  output     [7:0]    io_outputs_4_payload_1_0_2_6,
  output     [7:0]    io_outputs_4_payload_1_0_2_7,
  output     [7:0]    io_outputs_4_payload_1_0_2_8,
  output     [7:0]    io_outputs_4_payload_1_0_2_9,
  output     [7:0]    io_outputs_4_payload_1_0_2_10,
  output     [7:0]    io_outputs_4_payload_1_0_2_11,
  output     [7:0]    io_outputs_4_payload_1_0_2_12,
  output     [7:0]    io_outputs_4_payload_1_0_2_13,
  output     [7:0]    io_outputs_4_payload_1_0_2_14,
  output     [7:0]    io_outputs_4_payload_1_0_2_15,
  output     [7:0]    io_outputs_4_payload_1_1_0_0,
  output     [7:0]    io_outputs_4_payload_1_1_0_1,
  output     [7:0]    io_outputs_4_payload_1_1_0_2,
  output     [7:0]    io_outputs_4_payload_1_1_0_3,
  output     [7:0]    io_outputs_4_payload_1_1_0_4,
  output     [7:0]    io_outputs_4_payload_1_1_0_5,
  output     [7:0]    io_outputs_4_payload_1_1_0_6,
  output     [7:0]    io_outputs_4_payload_1_1_0_7,
  output     [7:0]    io_outputs_4_payload_1_1_0_8,
  output     [7:0]    io_outputs_4_payload_1_1_0_9,
  output     [7:0]    io_outputs_4_payload_1_1_0_10,
  output     [7:0]    io_outputs_4_payload_1_1_0_11,
  output     [7:0]    io_outputs_4_payload_1_1_0_12,
  output     [7:0]    io_outputs_4_payload_1_1_0_13,
  output     [7:0]    io_outputs_4_payload_1_1_0_14,
  output     [7:0]    io_outputs_4_payload_1_1_0_15,
  output     [7:0]    io_outputs_4_payload_1_1_1_0,
  output     [7:0]    io_outputs_4_payload_1_1_1_1,
  output     [7:0]    io_outputs_4_payload_1_1_1_2,
  output     [7:0]    io_outputs_4_payload_1_1_1_3,
  output     [7:0]    io_outputs_4_payload_1_1_1_4,
  output     [7:0]    io_outputs_4_payload_1_1_1_5,
  output     [7:0]    io_outputs_4_payload_1_1_1_6,
  output     [7:0]    io_outputs_4_payload_1_1_1_7,
  output     [7:0]    io_outputs_4_payload_1_1_1_8,
  output     [7:0]    io_outputs_4_payload_1_1_1_9,
  output     [7:0]    io_outputs_4_payload_1_1_1_10,
  output     [7:0]    io_outputs_4_payload_1_1_1_11,
  output     [7:0]    io_outputs_4_payload_1_1_1_12,
  output     [7:0]    io_outputs_4_payload_1_1_1_13,
  output     [7:0]    io_outputs_4_payload_1_1_1_14,
  output     [7:0]    io_outputs_4_payload_1_1_1_15,
  output     [7:0]    io_outputs_4_payload_1_1_2_0,
  output     [7:0]    io_outputs_4_payload_1_1_2_1,
  output     [7:0]    io_outputs_4_payload_1_1_2_2,
  output     [7:0]    io_outputs_4_payload_1_1_2_3,
  output     [7:0]    io_outputs_4_payload_1_1_2_4,
  output     [7:0]    io_outputs_4_payload_1_1_2_5,
  output     [7:0]    io_outputs_4_payload_1_1_2_6,
  output     [7:0]    io_outputs_4_payload_1_1_2_7,
  output     [7:0]    io_outputs_4_payload_1_1_2_8,
  output     [7:0]    io_outputs_4_payload_1_1_2_9,
  output     [7:0]    io_outputs_4_payload_1_1_2_10,
  output     [7:0]    io_outputs_4_payload_1_1_2_11,
  output     [7:0]    io_outputs_4_payload_1_1_2_12,
  output     [7:0]    io_outputs_4_payload_1_1_2_13,
  output     [7:0]    io_outputs_4_payload_1_1_2_14,
  output     [7:0]    io_outputs_4_payload_1_1_2_15,
  output     [7:0]    io_outputs_4_payload_1_2_0_0,
  output     [7:0]    io_outputs_4_payload_1_2_0_1,
  output     [7:0]    io_outputs_4_payload_1_2_0_2,
  output     [7:0]    io_outputs_4_payload_1_2_0_3,
  output     [7:0]    io_outputs_4_payload_1_2_0_4,
  output     [7:0]    io_outputs_4_payload_1_2_0_5,
  output     [7:0]    io_outputs_4_payload_1_2_0_6,
  output     [7:0]    io_outputs_4_payload_1_2_0_7,
  output     [7:0]    io_outputs_4_payload_1_2_0_8,
  output     [7:0]    io_outputs_4_payload_1_2_0_9,
  output     [7:0]    io_outputs_4_payload_1_2_0_10,
  output     [7:0]    io_outputs_4_payload_1_2_0_11,
  output     [7:0]    io_outputs_4_payload_1_2_0_12,
  output     [7:0]    io_outputs_4_payload_1_2_0_13,
  output     [7:0]    io_outputs_4_payload_1_2_0_14,
  output     [7:0]    io_outputs_4_payload_1_2_0_15,
  output     [7:0]    io_outputs_4_payload_1_2_1_0,
  output     [7:0]    io_outputs_4_payload_1_2_1_1,
  output     [7:0]    io_outputs_4_payload_1_2_1_2,
  output     [7:0]    io_outputs_4_payload_1_2_1_3,
  output     [7:0]    io_outputs_4_payload_1_2_1_4,
  output     [7:0]    io_outputs_4_payload_1_2_1_5,
  output     [7:0]    io_outputs_4_payload_1_2_1_6,
  output     [7:0]    io_outputs_4_payload_1_2_1_7,
  output     [7:0]    io_outputs_4_payload_1_2_1_8,
  output     [7:0]    io_outputs_4_payload_1_2_1_9,
  output     [7:0]    io_outputs_4_payload_1_2_1_10,
  output     [7:0]    io_outputs_4_payload_1_2_1_11,
  output     [7:0]    io_outputs_4_payload_1_2_1_12,
  output     [7:0]    io_outputs_4_payload_1_2_1_13,
  output     [7:0]    io_outputs_4_payload_1_2_1_14,
  output     [7:0]    io_outputs_4_payload_1_2_1_15,
  output     [7:0]    io_outputs_4_payload_1_2_2_0,
  output     [7:0]    io_outputs_4_payload_1_2_2_1,
  output     [7:0]    io_outputs_4_payload_1_2_2_2,
  output     [7:0]    io_outputs_4_payload_1_2_2_3,
  output     [7:0]    io_outputs_4_payload_1_2_2_4,
  output     [7:0]    io_outputs_4_payload_1_2_2_5,
  output     [7:0]    io_outputs_4_payload_1_2_2_6,
  output     [7:0]    io_outputs_4_payload_1_2_2_7,
  output     [7:0]    io_outputs_4_payload_1_2_2_8,
  output     [7:0]    io_outputs_4_payload_1_2_2_9,
  output     [7:0]    io_outputs_4_payload_1_2_2_10,
  output     [7:0]    io_outputs_4_payload_1_2_2_11,
  output     [7:0]    io_outputs_4_payload_1_2_2_12,
  output     [7:0]    io_outputs_4_payload_1_2_2_13,
  output     [7:0]    io_outputs_4_payload_1_2_2_14,
  output     [7:0]    io_outputs_4_payload_1_2_2_15,
  output reg          io_outputs_5_valid,
  input               io_outputs_5_ready,
  output     [7:0]    io_outputs_5_payload_0_0_0_0,
  output     [7:0]    io_outputs_5_payload_0_0_0_1,
  output     [7:0]    io_outputs_5_payload_0_0_0_2,
  output     [7:0]    io_outputs_5_payload_0_0_0_3,
  output     [7:0]    io_outputs_5_payload_0_0_0_4,
  output     [7:0]    io_outputs_5_payload_0_0_0_5,
  output     [7:0]    io_outputs_5_payload_0_0_0_6,
  output     [7:0]    io_outputs_5_payload_0_0_0_7,
  output     [7:0]    io_outputs_5_payload_0_0_0_8,
  output     [7:0]    io_outputs_5_payload_0_0_0_9,
  output     [7:0]    io_outputs_5_payload_0_0_0_10,
  output     [7:0]    io_outputs_5_payload_0_0_0_11,
  output     [7:0]    io_outputs_5_payload_0_0_0_12,
  output     [7:0]    io_outputs_5_payload_0_0_0_13,
  output     [7:0]    io_outputs_5_payload_0_0_0_14,
  output     [7:0]    io_outputs_5_payload_0_0_0_15,
  output     [7:0]    io_outputs_5_payload_0_0_1_0,
  output     [7:0]    io_outputs_5_payload_0_0_1_1,
  output     [7:0]    io_outputs_5_payload_0_0_1_2,
  output     [7:0]    io_outputs_5_payload_0_0_1_3,
  output     [7:0]    io_outputs_5_payload_0_0_1_4,
  output     [7:0]    io_outputs_5_payload_0_0_1_5,
  output     [7:0]    io_outputs_5_payload_0_0_1_6,
  output     [7:0]    io_outputs_5_payload_0_0_1_7,
  output     [7:0]    io_outputs_5_payload_0_0_1_8,
  output     [7:0]    io_outputs_5_payload_0_0_1_9,
  output     [7:0]    io_outputs_5_payload_0_0_1_10,
  output     [7:0]    io_outputs_5_payload_0_0_1_11,
  output     [7:0]    io_outputs_5_payload_0_0_1_12,
  output     [7:0]    io_outputs_5_payload_0_0_1_13,
  output     [7:0]    io_outputs_5_payload_0_0_1_14,
  output     [7:0]    io_outputs_5_payload_0_0_1_15,
  output     [7:0]    io_outputs_5_payload_0_0_2_0,
  output     [7:0]    io_outputs_5_payload_0_0_2_1,
  output     [7:0]    io_outputs_5_payload_0_0_2_2,
  output     [7:0]    io_outputs_5_payload_0_0_2_3,
  output     [7:0]    io_outputs_5_payload_0_0_2_4,
  output     [7:0]    io_outputs_5_payload_0_0_2_5,
  output     [7:0]    io_outputs_5_payload_0_0_2_6,
  output     [7:0]    io_outputs_5_payload_0_0_2_7,
  output     [7:0]    io_outputs_5_payload_0_0_2_8,
  output     [7:0]    io_outputs_5_payload_0_0_2_9,
  output     [7:0]    io_outputs_5_payload_0_0_2_10,
  output     [7:0]    io_outputs_5_payload_0_0_2_11,
  output     [7:0]    io_outputs_5_payload_0_0_2_12,
  output     [7:0]    io_outputs_5_payload_0_0_2_13,
  output     [7:0]    io_outputs_5_payload_0_0_2_14,
  output     [7:0]    io_outputs_5_payload_0_0_2_15,
  output     [7:0]    io_outputs_5_payload_0_1_0_0,
  output     [7:0]    io_outputs_5_payload_0_1_0_1,
  output     [7:0]    io_outputs_5_payload_0_1_0_2,
  output     [7:0]    io_outputs_5_payload_0_1_0_3,
  output     [7:0]    io_outputs_5_payload_0_1_0_4,
  output     [7:0]    io_outputs_5_payload_0_1_0_5,
  output     [7:0]    io_outputs_5_payload_0_1_0_6,
  output     [7:0]    io_outputs_5_payload_0_1_0_7,
  output     [7:0]    io_outputs_5_payload_0_1_0_8,
  output     [7:0]    io_outputs_5_payload_0_1_0_9,
  output     [7:0]    io_outputs_5_payload_0_1_0_10,
  output     [7:0]    io_outputs_5_payload_0_1_0_11,
  output     [7:0]    io_outputs_5_payload_0_1_0_12,
  output     [7:0]    io_outputs_5_payload_0_1_0_13,
  output     [7:0]    io_outputs_5_payload_0_1_0_14,
  output     [7:0]    io_outputs_5_payload_0_1_0_15,
  output     [7:0]    io_outputs_5_payload_0_1_1_0,
  output     [7:0]    io_outputs_5_payload_0_1_1_1,
  output     [7:0]    io_outputs_5_payload_0_1_1_2,
  output     [7:0]    io_outputs_5_payload_0_1_1_3,
  output     [7:0]    io_outputs_5_payload_0_1_1_4,
  output     [7:0]    io_outputs_5_payload_0_1_1_5,
  output     [7:0]    io_outputs_5_payload_0_1_1_6,
  output     [7:0]    io_outputs_5_payload_0_1_1_7,
  output     [7:0]    io_outputs_5_payload_0_1_1_8,
  output     [7:0]    io_outputs_5_payload_0_1_1_9,
  output     [7:0]    io_outputs_5_payload_0_1_1_10,
  output     [7:0]    io_outputs_5_payload_0_1_1_11,
  output     [7:0]    io_outputs_5_payload_0_1_1_12,
  output     [7:0]    io_outputs_5_payload_0_1_1_13,
  output     [7:0]    io_outputs_5_payload_0_1_1_14,
  output     [7:0]    io_outputs_5_payload_0_1_1_15,
  output     [7:0]    io_outputs_5_payload_0_1_2_0,
  output     [7:0]    io_outputs_5_payload_0_1_2_1,
  output     [7:0]    io_outputs_5_payload_0_1_2_2,
  output     [7:0]    io_outputs_5_payload_0_1_2_3,
  output     [7:0]    io_outputs_5_payload_0_1_2_4,
  output     [7:0]    io_outputs_5_payload_0_1_2_5,
  output     [7:0]    io_outputs_5_payload_0_1_2_6,
  output     [7:0]    io_outputs_5_payload_0_1_2_7,
  output     [7:0]    io_outputs_5_payload_0_1_2_8,
  output     [7:0]    io_outputs_5_payload_0_1_2_9,
  output     [7:0]    io_outputs_5_payload_0_1_2_10,
  output     [7:0]    io_outputs_5_payload_0_1_2_11,
  output     [7:0]    io_outputs_5_payload_0_1_2_12,
  output     [7:0]    io_outputs_5_payload_0_1_2_13,
  output     [7:0]    io_outputs_5_payload_0_1_2_14,
  output     [7:0]    io_outputs_5_payload_0_1_2_15,
  output     [7:0]    io_outputs_5_payload_0_2_0_0,
  output     [7:0]    io_outputs_5_payload_0_2_0_1,
  output     [7:0]    io_outputs_5_payload_0_2_0_2,
  output     [7:0]    io_outputs_5_payload_0_2_0_3,
  output     [7:0]    io_outputs_5_payload_0_2_0_4,
  output     [7:0]    io_outputs_5_payload_0_2_0_5,
  output     [7:0]    io_outputs_5_payload_0_2_0_6,
  output     [7:0]    io_outputs_5_payload_0_2_0_7,
  output     [7:0]    io_outputs_5_payload_0_2_0_8,
  output     [7:0]    io_outputs_5_payload_0_2_0_9,
  output     [7:0]    io_outputs_5_payload_0_2_0_10,
  output     [7:0]    io_outputs_5_payload_0_2_0_11,
  output     [7:0]    io_outputs_5_payload_0_2_0_12,
  output     [7:0]    io_outputs_5_payload_0_2_0_13,
  output     [7:0]    io_outputs_5_payload_0_2_0_14,
  output     [7:0]    io_outputs_5_payload_0_2_0_15,
  output     [7:0]    io_outputs_5_payload_0_2_1_0,
  output     [7:0]    io_outputs_5_payload_0_2_1_1,
  output     [7:0]    io_outputs_5_payload_0_2_1_2,
  output     [7:0]    io_outputs_5_payload_0_2_1_3,
  output     [7:0]    io_outputs_5_payload_0_2_1_4,
  output     [7:0]    io_outputs_5_payload_0_2_1_5,
  output     [7:0]    io_outputs_5_payload_0_2_1_6,
  output     [7:0]    io_outputs_5_payload_0_2_1_7,
  output     [7:0]    io_outputs_5_payload_0_2_1_8,
  output     [7:0]    io_outputs_5_payload_0_2_1_9,
  output     [7:0]    io_outputs_5_payload_0_2_1_10,
  output     [7:0]    io_outputs_5_payload_0_2_1_11,
  output     [7:0]    io_outputs_5_payload_0_2_1_12,
  output     [7:0]    io_outputs_5_payload_0_2_1_13,
  output     [7:0]    io_outputs_5_payload_0_2_1_14,
  output     [7:0]    io_outputs_5_payload_0_2_1_15,
  output     [7:0]    io_outputs_5_payload_0_2_2_0,
  output     [7:0]    io_outputs_5_payload_0_2_2_1,
  output     [7:0]    io_outputs_5_payload_0_2_2_2,
  output     [7:0]    io_outputs_5_payload_0_2_2_3,
  output     [7:0]    io_outputs_5_payload_0_2_2_4,
  output     [7:0]    io_outputs_5_payload_0_2_2_5,
  output     [7:0]    io_outputs_5_payload_0_2_2_6,
  output     [7:0]    io_outputs_5_payload_0_2_2_7,
  output     [7:0]    io_outputs_5_payload_0_2_2_8,
  output     [7:0]    io_outputs_5_payload_0_2_2_9,
  output     [7:0]    io_outputs_5_payload_0_2_2_10,
  output     [7:0]    io_outputs_5_payload_0_2_2_11,
  output     [7:0]    io_outputs_5_payload_0_2_2_12,
  output     [7:0]    io_outputs_5_payload_0_2_2_13,
  output     [7:0]    io_outputs_5_payload_0_2_2_14,
  output     [7:0]    io_outputs_5_payload_0_2_2_15,
  output     [7:0]    io_outputs_5_payload_1_0_0_0,
  output     [7:0]    io_outputs_5_payload_1_0_0_1,
  output     [7:0]    io_outputs_5_payload_1_0_0_2,
  output     [7:0]    io_outputs_5_payload_1_0_0_3,
  output     [7:0]    io_outputs_5_payload_1_0_0_4,
  output     [7:0]    io_outputs_5_payload_1_0_0_5,
  output     [7:0]    io_outputs_5_payload_1_0_0_6,
  output     [7:0]    io_outputs_5_payload_1_0_0_7,
  output     [7:0]    io_outputs_5_payload_1_0_0_8,
  output     [7:0]    io_outputs_5_payload_1_0_0_9,
  output     [7:0]    io_outputs_5_payload_1_0_0_10,
  output     [7:0]    io_outputs_5_payload_1_0_0_11,
  output     [7:0]    io_outputs_5_payload_1_0_0_12,
  output     [7:0]    io_outputs_5_payload_1_0_0_13,
  output     [7:0]    io_outputs_5_payload_1_0_0_14,
  output     [7:0]    io_outputs_5_payload_1_0_0_15,
  output     [7:0]    io_outputs_5_payload_1_0_1_0,
  output     [7:0]    io_outputs_5_payload_1_0_1_1,
  output     [7:0]    io_outputs_5_payload_1_0_1_2,
  output     [7:0]    io_outputs_5_payload_1_0_1_3,
  output     [7:0]    io_outputs_5_payload_1_0_1_4,
  output     [7:0]    io_outputs_5_payload_1_0_1_5,
  output     [7:0]    io_outputs_5_payload_1_0_1_6,
  output     [7:0]    io_outputs_5_payload_1_0_1_7,
  output     [7:0]    io_outputs_5_payload_1_0_1_8,
  output     [7:0]    io_outputs_5_payload_1_0_1_9,
  output     [7:0]    io_outputs_5_payload_1_0_1_10,
  output     [7:0]    io_outputs_5_payload_1_0_1_11,
  output     [7:0]    io_outputs_5_payload_1_0_1_12,
  output     [7:0]    io_outputs_5_payload_1_0_1_13,
  output     [7:0]    io_outputs_5_payload_1_0_1_14,
  output     [7:0]    io_outputs_5_payload_1_0_1_15,
  output     [7:0]    io_outputs_5_payload_1_0_2_0,
  output     [7:0]    io_outputs_5_payload_1_0_2_1,
  output     [7:0]    io_outputs_5_payload_1_0_2_2,
  output     [7:0]    io_outputs_5_payload_1_0_2_3,
  output     [7:0]    io_outputs_5_payload_1_0_2_4,
  output     [7:0]    io_outputs_5_payload_1_0_2_5,
  output     [7:0]    io_outputs_5_payload_1_0_2_6,
  output     [7:0]    io_outputs_5_payload_1_0_2_7,
  output     [7:0]    io_outputs_5_payload_1_0_2_8,
  output     [7:0]    io_outputs_5_payload_1_0_2_9,
  output     [7:0]    io_outputs_5_payload_1_0_2_10,
  output     [7:0]    io_outputs_5_payload_1_0_2_11,
  output     [7:0]    io_outputs_5_payload_1_0_2_12,
  output     [7:0]    io_outputs_5_payload_1_0_2_13,
  output     [7:0]    io_outputs_5_payload_1_0_2_14,
  output     [7:0]    io_outputs_5_payload_1_0_2_15,
  output     [7:0]    io_outputs_5_payload_1_1_0_0,
  output     [7:0]    io_outputs_5_payload_1_1_0_1,
  output     [7:0]    io_outputs_5_payload_1_1_0_2,
  output     [7:0]    io_outputs_5_payload_1_1_0_3,
  output     [7:0]    io_outputs_5_payload_1_1_0_4,
  output     [7:0]    io_outputs_5_payload_1_1_0_5,
  output     [7:0]    io_outputs_5_payload_1_1_0_6,
  output     [7:0]    io_outputs_5_payload_1_1_0_7,
  output     [7:0]    io_outputs_5_payload_1_1_0_8,
  output     [7:0]    io_outputs_5_payload_1_1_0_9,
  output     [7:0]    io_outputs_5_payload_1_1_0_10,
  output     [7:0]    io_outputs_5_payload_1_1_0_11,
  output     [7:0]    io_outputs_5_payload_1_1_0_12,
  output     [7:0]    io_outputs_5_payload_1_1_0_13,
  output     [7:0]    io_outputs_5_payload_1_1_0_14,
  output     [7:0]    io_outputs_5_payload_1_1_0_15,
  output     [7:0]    io_outputs_5_payload_1_1_1_0,
  output     [7:0]    io_outputs_5_payload_1_1_1_1,
  output     [7:0]    io_outputs_5_payload_1_1_1_2,
  output     [7:0]    io_outputs_5_payload_1_1_1_3,
  output     [7:0]    io_outputs_5_payload_1_1_1_4,
  output     [7:0]    io_outputs_5_payload_1_1_1_5,
  output     [7:0]    io_outputs_5_payload_1_1_1_6,
  output     [7:0]    io_outputs_5_payload_1_1_1_7,
  output     [7:0]    io_outputs_5_payload_1_1_1_8,
  output     [7:0]    io_outputs_5_payload_1_1_1_9,
  output     [7:0]    io_outputs_5_payload_1_1_1_10,
  output     [7:0]    io_outputs_5_payload_1_1_1_11,
  output     [7:0]    io_outputs_5_payload_1_1_1_12,
  output     [7:0]    io_outputs_5_payload_1_1_1_13,
  output     [7:0]    io_outputs_5_payload_1_1_1_14,
  output     [7:0]    io_outputs_5_payload_1_1_1_15,
  output     [7:0]    io_outputs_5_payload_1_1_2_0,
  output     [7:0]    io_outputs_5_payload_1_1_2_1,
  output     [7:0]    io_outputs_5_payload_1_1_2_2,
  output     [7:0]    io_outputs_5_payload_1_1_2_3,
  output     [7:0]    io_outputs_5_payload_1_1_2_4,
  output     [7:0]    io_outputs_5_payload_1_1_2_5,
  output     [7:0]    io_outputs_5_payload_1_1_2_6,
  output     [7:0]    io_outputs_5_payload_1_1_2_7,
  output     [7:0]    io_outputs_5_payload_1_1_2_8,
  output     [7:0]    io_outputs_5_payload_1_1_2_9,
  output     [7:0]    io_outputs_5_payload_1_1_2_10,
  output     [7:0]    io_outputs_5_payload_1_1_2_11,
  output     [7:0]    io_outputs_5_payload_1_1_2_12,
  output     [7:0]    io_outputs_5_payload_1_1_2_13,
  output     [7:0]    io_outputs_5_payload_1_1_2_14,
  output     [7:0]    io_outputs_5_payload_1_1_2_15,
  output     [7:0]    io_outputs_5_payload_1_2_0_0,
  output     [7:0]    io_outputs_5_payload_1_2_0_1,
  output     [7:0]    io_outputs_5_payload_1_2_0_2,
  output     [7:0]    io_outputs_5_payload_1_2_0_3,
  output     [7:0]    io_outputs_5_payload_1_2_0_4,
  output     [7:0]    io_outputs_5_payload_1_2_0_5,
  output     [7:0]    io_outputs_5_payload_1_2_0_6,
  output     [7:0]    io_outputs_5_payload_1_2_0_7,
  output     [7:0]    io_outputs_5_payload_1_2_0_8,
  output     [7:0]    io_outputs_5_payload_1_2_0_9,
  output     [7:0]    io_outputs_5_payload_1_2_0_10,
  output     [7:0]    io_outputs_5_payload_1_2_0_11,
  output     [7:0]    io_outputs_5_payload_1_2_0_12,
  output     [7:0]    io_outputs_5_payload_1_2_0_13,
  output     [7:0]    io_outputs_5_payload_1_2_0_14,
  output     [7:0]    io_outputs_5_payload_1_2_0_15,
  output     [7:0]    io_outputs_5_payload_1_2_1_0,
  output     [7:0]    io_outputs_5_payload_1_2_1_1,
  output     [7:0]    io_outputs_5_payload_1_2_1_2,
  output     [7:0]    io_outputs_5_payload_1_2_1_3,
  output     [7:0]    io_outputs_5_payload_1_2_1_4,
  output     [7:0]    io_outputs_5_payload_1_2_1_5,
  output     [7:0]    io_outputs_5_payload_1_2_1_6,
  output     [7:0]    io_outputs_5_payload_1_2_1_7,
  output     [7:0]    io_outputs_5_payload_1_2_1_8,
  output     [7:0]    io_outputs_5_payload_1_2_1_9,
  output     [7:0]    io_outputs_5_payload_1_2_1_10,
  output     [7:0]    io_outputs_5_payload_1_2_1_11,
  output     [7:0]    io_outputs_5_payload_1_2_1_12,
  output     [7:0]    io_outputs_5_payload_1_2_1_13,
  output     [7:0]    io_outputs_5_payload_1_2_1_14,
  output     [7:0]    io_outputs_5_payload_1_2_1_15,
  output     [7:0]    io_outputs_5_payload_1_2_2_0,
  output     [7:0]    io_outputs_5_payload_1_2_2_1,
  output     [7:0]    io_outputs_5_payload_1_2_2_2,
  output     [7:0]    io_outputs_5_payload_1_2_2_3,
  output     [7:0]    io_outputs_5_payload_1_2_2_4,
  output     [7:0]    io_outputs_5_payload_1_2_2_5,
  output     [7:0]    io_outputs_5_payload_1_2_2_6,
  output     [7:0]    io_outputs_5_payload_1_2_2_7,
  output     [7:0]    io_outputs_5_payload_1_2_2_8,
  output     [7:0]    io_outputs_5_payload_1_2_2_9,
  output     [7:0]    io_outputs_5_payload_1_2_2_10,
  output     [7:0]    io_outputs_5_payload_1_2_2_11,
  output     [7:0]    io_outputs_5_payload_1_2_2_12,
  output     [7:0]    io_outputs_5_payload_1_2_2_13,
  output     [7:0]    io_outputs_5_payload_1_2_2_14,
  output     [7:0]    io_outputs_5_payload_1_2_2_15,
  output reg          io_outputs_6_valid,
  input               io_outputs_6_ready,
  output     [7:0]    io_outputs_6_payload_0_0_0_0,
  output     [7:0]    io_outputs_6_payload_0_0_0_1,
  output     [7:0]    io_outputs_6_payload_0_0_0_2,
  output     [7:0]    io_outputs_6_payload_0_0_0_3,
  output     [7:0]    io_outputs_6_payload_0_0_0_4,
  output     [7:0]    io_outputs_6_payload_0_0_0_5,
  output     [7:0]    io_outputs_6_payload_0_0_0_6,
  output     [7:0]    io_outputs_6_payload_0_0_0_7,
  output     [7:0]    io_outputs_6_payload_0_0_0_8,
  output     [7:0]    io_outputs_6_payload_0_0_0_9,
  output     [7:0]    io_outputs_6_payload_0_0_0_10,
  output     [7:0]    io_outputs_6_payload_0_0_0_11,
  output     [7:0]    io_outputs_6_payload_0_0_0_12,
  output     [7:0]    io_outputs_6_payload_0_0_0_13,
  output     [7:0]    io_outputs_6_payload_0_0_0_14,
  output     [7:0]    io_outputs_6_payload_0_0_0_15,
  output     [7:0]    io_outputs_6_payload_0_0_1_0,
  output     [7:0]    io_outputs_6_payload_0_0_1_1,
  output     [7:0]    io_outputs_6_payload_0_0_1_2,
  output     [7:0]    io_outputs_6_payload_0_0_1_3,
  output     [7:0]    io_outputs_6_payload_0_0_1_4,
  output     [7:0]    io_outputs_6_payload_0_0_1_5,
  output     [7:0]    io_outputs_6_payload_0_0_1_6,
  output     [7:0]    io_outputs_6_payload_0_0_1_7,
  output     [7:0]    io_outputs_6_payload_0_0_1_8,
  output     [7:0]    io_outputs_6_payload_0_0_1_9,
  output     [7:0]    io_outputs_6_payload_0_0_1_10,
  output     [7:0]    io_outputs_6_payload_0_0_1_11,
  output     [7:0]    io_outputs_6_payload_0_0_1_12,
  output     [7:0]    io_outputs_6_payload_0_0_1_13,
  output     [7:0]    io_outputs_6_payload_0_0_1_14,
  output     [7:0]    io_outputs_6_payload_0_0_1_15,
  output     [7:0]    io_outputs_6_payload_0_0_2_0,
  output     [7:0]    io_outputs_6_payload_0_0_2_1,
  output     [7:0]    io_outputs_6_payload_0_0_2_2,
  output     [7:0]    io_outputs_6_payload_0_0_2_3,
  output     [7:0]    io_outputs_6_payload_0_0_2_4,
  output     [7:0]    io_outputs_6_payload_0_0_2_5,
  output     [7:0]    io_outputs_6_payload_0_0_2_6,
  output     [7:0]    io_outputs_6_payload_0_0_2_7,
  output     [7:0]    io_outputs_6_payload_0_0_2_8,
  output     [7:0]    io_outputs_6_payload_0_0_2_9,
  output     [7:0]    io_outputs_6_payload_0_0_2_10,
  output     [7:0]    io_outputs_6_payload_0_0_2_11,
  output     [7:0]    io_outputs_6_payload_0_0_2_12,
  output     [7:0]    io_outputs_6_payload_0_0_2_13,
  output     [7:0]    io_outputs_6_payload_0_0_2_14,
  output     [7:0]    io_outputs_6_payload_0_0_2_15,
  output     [7:0]    io_outputs_6_payload_0_1_0_0,
  output     [7:0]    io_outputs_6_payload_0_1_0_1,
  output     [7:0]    io_outputs_6_payload_0_1_0_2,
  output     [7:0]    io_outputs_6_payload_0_1_0_3,
  output     [7:0]    io_outputs_6_payload_0_1_0_4,
  output     [7:0]    io_outputs_6_payload_0_1_0_5,
  output     [7:0]    io_outputs_6_payload_0_1_0_6,
  output     [7:0]    io_outputs_6_payload_0_1_0_7,
  output     [7:0]    io_outputs_6_payload_0_1_0_8,
  output     [7:0]    io_outputs_6_payload_0_1_0_9,
  output     [7:0]    io_outputs_6_payload_0_1_0_10,
  output     [7:0]    io_outputs_6_payload_0_1_0_11,
  output     [7:0]    io_outputs_6_payload_0_1_0_12,
  output     [7:0]    io_outputs_6_payload_0_1_0_13,
  output     [7:0]    io_outputs_6_payload_0_1_0_14,
  output     [7:0]    io_outputs_6_payload_0_1_0_15,
  output     [7:0]    io_outputs_6_payload_0_1_1_0,
  output     [7:0]    io_outputs_6_payload_0_1_1_1,
  output     [7:0]    io_outputs_6_payload_0_1_1_2,
  output     [7:0]    io_outputs_6_payload_0_1_1_3,
  output     [7:0]    io_outputs_6_payload_0_1_1_4,
  output     [7:0]    io_outputs_6_payload_0_1_1_5,
  output     [7:0]    io_outputs_6_payload_0_1_1_6,
  output     [7:0]    io_outputs_6_payload_0_1_1_7,
  output     [7:0]    io_outputs_6_payload_0_1_1_8,
  output     [7:0]    io_outputs_6_payload_0_1_1_9,
  output     [7:0]    io_outputs_6_payload_0_1_1_10,
  output     [7:0]    io_outputs_6_payload_0_1_1_11,
  output     [7:0]    io_outputs_6_payload_0_1_1_12,
  output     [7:0]    io_outputs_6_payload_0_1_1_13,
  output     [7:0]    io_outputs_6_payload_0_1_1_14,
  output     [7:0]    io_outputs_6_payload_0_1_1_15,
  output     [7:0]    io_outputs_6_payload_0_1_2_0,
  output     [7:0]    io_outputs_6_payload_0_1_2_1,
  output     [7:0]    io_outputs_6_payload_0_1_2_2,
  output     [7:0]    io_outputs_6_payload_0_1_2_3,
  output     [7:0]    io_outputs_6_payload_0_1_2_4,
  output     [7:0]    io_outputs_6_payload_0_1_2_5,
  output     [7:0]    io_outputs_6_payload_0_1_2_6,
  output     [7:0]    io_outputs_6_payload_0_1_2_7,
  output     [7:0]    io_outputs_6_payload_0_1_2_8,
  output     [7:0]    io_outputs_6_payload_0_1_2_9,
  output     [7:0]    io_outputs_6_payload_0_1_2_10,
  output     [7:0]    io_outputs_6_payload_0_1_2_11,
  output     [7:0]    io_outputs_6_payload_0_1_2_12,
  output     [7:0]    io_outputs_6_payload_0_1_2_13,
  output     [7:0]    io_outputs_6_payload_0_1_2_14,
  output     [7:0]    io_outputs_6_payload_0_1_2_15,
  output     [7:0]    io_outputs_6_payload_0_2_0_0,
  output     [7:0]    io_outputs_6_payload_0_2_0_1,
  output     [7:0]    io_outputs_6_payload_0_2_0_2,
  output     [7:0]    io_outputs_6_payload_0_2_0_3,
  output     [7:0]    io_outputs_6_payload_0_2_0_4,
  output     [7:0]    io_outputs_6_payload_0_2_0_5,
  output     [7:0]    io_outputs_6_payload_0_2_0_6,
  output     [7:0]    io_outputs_6_payload_0_2_0_7,
  output     [7:0]    io_outputs_6_payload_0_2_0_8,
  output     [7:0]    io_outputs_6_payload_0_2_0_9,
  output     [7:0]    io_outputs_6_payload_0_2_0_10,
  output     [7:0]    io_outputs_6_payload_0_2_0_11,
  output     [7:0]    io_outputs_6_payload_0_2_0_12,
  output     [7:0]    io_outputs_6_payload_0_2_0_13,
  output     [7:0]    io_outputs_6_payload_0_2_0_14,
  output     [7:0]    io_outputs_6_payload_0_2_0_15,
  output     [7:0]    io_outputs_6_payload_0_2_1_0,
  output     [7:0]    io_outputs_6_payload_0_2_1_1,
  output     [7:0]    io_outputs_6_payload_0_2_1_2,
  output     [7:0]    io_outputs_6_payload_0_2_1_3,
  output     [7:0]    io_outputs_6_payload_0_2_1_4,
  output     [7:0]    io_outputs_6_payload_0_2_1_5,
  output     [7:0]    io_outputs_6_payload_0_2_1_6,
  output     [7:0]    io_outputs_6_payload_0_2_1_7,
  output     [7:0]    io_outputs_6_payload_0_2_1_8,
  output     [7:0]    io_outputs_6_payload_0_2_1_9,
  output     [7:0]    io_outputs_6_payload_0_2_1_10,
  output     [7:0]    io_outputs_6_payload_0_2_1_11,
  output     [7:0]    io_outputs_6_payload_0_2_1_12,
  output     [7:0]    io_outputs_6_payload_0_2_1_13,
  output     [7:0]    io_outputs_6_payload_0_2_1_14,
  output     [7:0]    io_outputs_6_payload_0_2_1_15,
  output     [7:0]    io_outputs_6_payload_0_2_2_0,
  output     [7:0]    io_outputs_6_payload_0_2_2_1,
  output     [7:0]    io_outputs_6_payload_0_2_2_2,
  output     [7:0]    io_outputs_6_payload_0_2_2_3,
  output     [7:0]    io_outputs_6_payload_0_2_2_4,
  output     [7:0]    io_outputs_6_payload_0_2_2_5,
  output     [7:0]    io_outputs_6_payload_0_2_2_6,
  output     [7:0]    io_outputs_6_payload_0_2_2_7,
  output     [7:0]    io_outputs_6_payload_0_2_2_8,
  output     [7:0]    io_outputs_6_payload_0_2_2_9,
  output     [7:0]    io_outputs_6_payload_0_2_2_10,
  output     [7:0]    io_outputs_6_payload_0_2_2_11,
  output     [7:0]    io_outputs_6_payload_0_2_2_12,
  output     [7:0]    io_outputs_6_payload_0_2_2_13,
  output     [7:0]    io_outputs_6_payload_0_2_2_14,
  output     [7:0]    io_outputs_6_payload_0_2_2_15,
  output     [7:0]    io_outputs_6_payload_1_0_0_0,
  output     [7:0]    io_outputs_6_payload_1_0_0_1,
  output     [7:0]    io_outputs_6_payload_1_0_0_2,
  output     [7:0]    io_outputs_6_payload_1_0_0_3,
  output     [7:0]    io_outputs_6_payload_1_0_0_4,
  output     [7:0]    io_outputs_6_payload_1_0_0_5,
  output     [7:0]    io_outputs_6_payload_1_0_0_6,
  output     [7:0]    io_outputs_6_payload_1_0_0_7,
  output     [7:0]    io_outputs_6_payload_1_0_0_8,
  output     [7:0]    io_outputs_6_payload_1_0_0_9,
  output     [7:0]    io_outputs_6_payload_1_0_0_10,
  output     [7:0]    io_outputs_6_payload_1_0_0_11,
  output     [7:0]    io_outputs_6_payload_1_0_0_12,
  output     [7:0]    io_outputs_6_payload_1_0_0_13,
  output     [7:0]    io_outputs_6_payload_1_0_0_14,
  output     [7:0]    io_outputs_6_payload_1_0_0_15,
  output     [7:0]    io_outputs_6_payload_1_0_1_0,
  output     [7:0]    io_outputs_6_payload_1_0_1_1,
  output     [7:0]    io_outputs_6_payload_1_0_1_2,
  output     [7:0]    io_outputs_6_payload_1_0_1_3,
  output     [7:0]    io_outputs_6_payload_1_0_1_4,
  output     [7:0]    io_outputs_6_payload_1_0_1_5,
  output     [7:0]    io_outputs_6_payload_1_0_1_6,
  output     [7:0]    io_outputs_6_payload_1_0_1_7,
  output     [7:0]    io_outputs_6_payload_1_0_1_8,
  output     [7:0]    io_outputs_6_payload_1_0_1_9,
  output     [7:0]    io_outputs_6_payload_1_0_1_10,
  output     [7:0]    io_outputs_6_payload_1_0_1_11,
  output     [7:0]    io_outputs_6_payload_1_0_1_12,
  output     [7:0]    io_outputs_6_payload_1_0_1_13,
  output     [7:0]    io_outputs_6_payload_1_0_1_14,
  output     [7:0]    io_outputs_6_payload_1_0_1_15,
  output     [7:0]    io_outputs_6_payload_1_0_2_0,
  output     [7:0]    io_outputs_6_payload_1_0_2_1,
  output     [7:0]    io_outputs_6_payload_1_0_2_2,
  output     [7:0]    io_outputs_6_payload_1_0_2_3,
  output     [7:0]    io_outputs_6_payload_1_0_2_4,
  output     [7:0]    io_outputs_6_payload_1_0_2_5,
  output     [7:0]    io_outputs_6_payload_1_0_2_6,
  output     [7:0]    io_outputs_6_payload_1_0_2_7,
  output     [7:0]    io_outputs_6_payload_1_0_2_8,
  output     [7:0]    io_outputs_6_payload_1_0_2_9,
  output     [7:0]    io_outputs_6_payload_1_0_2_10,
  output     [7:0]    io_outputs_6_payload_1_0_2_11,
  output     [7:0]    io_outputs_6_payload_1_0_2_12,
  output     [7:0]    io_outputs_6_payload_1_0_2_13,
  output     [7:0]    io_outputs_6_payload_1_0_2_14,
  output     [7:0]    io_outputs_6_payload_1_0_2_15,
  output     [7:0]    io_outputs_6_payload_1_1_0_0,
  output     [7:0]    io_outputs_6_payload_1_1_0_1,
  output     [7:0]    io_outputs_6_payload_1_1_0_2,
  output     [7:0]    io_outputs_6_payload_1_1_0_3,
  output     [7:0]    io_outputs_6_payload_1_1_0_4,
  output     [7:0]    io_outputs_6_payload_1_1_0_5,
  output     [7:0]    io_outputs_6_payload_1_1_0_6,
  output     [7:0]    io_outputs_6_payload_1_1_0_7,
  output     [7:0]    io_outputs_6_payload_1_1_0_8,
  output     [7:0]    io_outputs_6_payload_1_1_0_9,
  output     [7:0]    io_outputs_6_payload_1_1_0_10,
  output     [7:0]    io_outputs_6_payload_1_1_0_11,
  output     [7:0]    io_outputs_6_payload_1_1_0_12,
  output     [7:0]    io_outputs_6_payload_1_1_0_13,
  output     [7:0]    io_outputs_6_payload_1_1_0_14,
  output     [7:0]    io_outputs_6_payload_1_1_0_15,
  output     [7:0]    io_outputs_6_payload_1_1_1_0,
  output     [7:0]    io_outputs_6_payload_1_1_1_1,
  output     [7:0]    io_outputs_6_payload_1_1_1_2,
  output     [7:0]    io_outputs_6_payload_1_1_1_3,
  output     [7:0]    io_outputs_6_payload_1_1_1_4,
  output     [7:0]    io_outputs_6_payload_1_1_1_5,
  output     [7:0]    io_outputs_6_payload_1_1_1_6,
  output     [7:0]    io_outputs_6_payload_1_1_1_7,
  output     [7:0]    io_outputs_6_payload_1_1_1_8,
  output     [7:0]    io_outputs_6_payload_1_1_1_9,
  output     [7:0]    io_outputs_6_payload_1_1_1_10,
  output     [7:0]    io_outputs_6_payload_1_1_1_11,
  output     [7:0]    io_outputs_6_payload_1_1_1_12,
  output     [7:0]    io_outputs_6_payload_1_1_1_13,
  output     [7:0]    io_outputs_6_payload_1_1_1_14,
  output     [7:0]    io_outputs_6_payload_1_1_1_15,
  output     [7:0]    io_outputs_6_payload_1_1_2_0,
  output     [7:0]    io_outputs_6_payload_1_1_2_1,
  output     [7:0]    io_outputs_6_payload_1_1_2_2,
  output     [7:0]    io_outputs_6_payload_1_1_2_3,
  output     [7:0]    io_outputs_6_payload_1_1_2_4,
  output     [7:0]    io_outputs_6_payload_1_1_2_5,
  output     [7:0]    io_outputs_6_payload_1_1_2_6,
  output     [7:0]    io_outputs_6_payload_1_1_2_7,
  output     [7:0]    io_outputs_6_payload_1_1_2_8,
  output     [7:0]    io_outputs_6_payload_1_1_2_9,
  output     [7:0]    io_outputs_6_payload_1_1_2_10,
  output     [7:0]    io_outputs_6_payload_1_1_2_11,
  output     [7:0]    io_outputs_6_payload_1_1_2_12,
  output     [7:0]    io_outputs_6_payload_1_1_2_13,
  output     [7:0]    io_outputs_6_payload_1_1_2_14,
  output     [7:0]    io_outputs_6_payload_1_1_2_15,
  output     [7:0]    io_outputs_6_payload_1_2_0_0,
  output     [7:0]    io_outputs_6_payload_1_2_0_1,
  output     [7:0]    io_outputs_6_payload_1_2_0_2,
  output     [7:0]    io_outputs_6_payload_1_2_0_3,
  output     [7:0]    io_outputs_6_payload_1_2_0_4,
  output     [7:0]    io_outputs_6_payload_1_2_0_5,
  output     [7:0]    io_outputs_6_payload_1_2_0_6,
  output     [7:0]    io_outputs_6_payload_1_2_0_7,
  output     [7:0]    io_outputs_6_payload_1_2_0_8,
  output     [7:0]    io_outputs_6_payload_1_2_0_9,
  output     [7:0]    io_outputs_6_payload_1_2_0_10,
  output     [7:0]    io_outputs_6_payload_1_2_0_11,
  output     [7:0]    io_outputs_6_payload_1_2_0_12,
  output     [7:0]    io_outputs_6_payload_1_2_0_13,
  output     [7:0]    io_outputs_6_payload_1_2_0_14,
  output     [7:0]    io_outputs_6_payload_1_2_0_15,
  output     [7:0]    io_outputs_6_payload_1_2_1_0,
  output     [7:0]    io_outputs_6_payload_1_2_1_1,
  output     [7:0]    io_outputs_6_payload_1_2_1_2,
  output     [7:0]    io_outputs_6_payload_1_2_1_3,
  output     [7:0]    io_outputs_6_payload_1_2_1_4,
  output     [7:0]    io_outputs_6_payload_1_2_1_5,
  output     [7:0]    io_outputs_6_payload_1_2_1_6,
  output     [7:0]    io_outputs_6_payload_1_2_1_7,
  output     [7:0]    io_outputs_6_payload_1_2_1_8,
  output     [7:0]    io_outputs_6_payload_1_2_1_9,
  output     [7:0]    io_outputs_6_payload_1_2_1_10,
  output     [7:0]    io_outputs_6_payload_1_2_1_11,
  output     [7:0]    io_outputs_6_payload_1_2_1_12,
  output     [7:0]    io_outputs_6_payload_1_2_1_13,
  output     [7:0]    io_outputs_6_payload_1_2_1_14,
  output     [7:0]    io_outputs_6_payload_1_2_1_15,
  output     [7:0]    io_outputs_6_payload_1_2_2_0,
  output     [7:0]    io_outputs_6_payload_1_2_2_1,
  output     [7:0]    io_outputs_6_payload_1_2_2_2,
  output     [7:0]    io_outputs_6_payload_1_2_2_3,
  output     [7:0]    io_outputs_6_payload_1_2_2_4,
  output     [7:0]    io_outputs_6_payload_1_2_2_5,
  output     [7:0]    io_outputs_6_payload_1_2_2_6,
  output     [7:0]    io_outputs_6_payload_1_2_2_7,
  output     [7:0]    io_outputs_6_payload_1_2_2_8,
  output     [7:0]    io_outputs_6_payload_1_2_2_9,
  output     [7:0]    io_outputs_6_payload_1_2_2_10,
  output     [7:0]    io_outputs_6_payload_1_2_2_11,
  output     [7:0]    io_outputs_6_payload_1_2_2_12,
  output     [7:0]    io_outputs_6_payload_1_2_2_13,
  output     [7:0]    io_outputs_6_payload_1_2_2_14,
  output     [7:0]    io_outputs_6_payload_1_2_2_15,
  output reg          io_outputs_7_valid,
  input               io_outputs_7_ready,
  output     [7:0]    io_outputs_7_payload_0_0_0_0,
  output     [7:0]    io_outputs_7_payload_0_0_0_1,
  output     [7:0]    io_outputs_7_payload_0_0_0_2,
  output     [7:0]    io_outputs_7_payload_0_0_0_3,
  output     [7:0]    io_outputs_7_payload_0_0_0_4,
  output     [7:0]    io_outputs_7_payload_0_0_0_5,
  output     [7:0]    io_outputs_7_payload_0_0_0_6,
  output     [7:0]    io_outputs_7_payload_0_0_0_7,
  output     [7:0]    io_outputs_7_payload_0_0_0_8,
  output     [7:0]    io_outputs_7_payload_0_0_0_9,
  output     [7:0]    io_outputs_7_payload_0_0_0_10,
  output     [7:0]    io_outputs_7_payload_0_0_0_11,
  output     [7:0]    io_outputs_7_payload_0_0_0_12,
  output     [7:0]    io_outputs_7_payload_0_0_0_13,
  output     [7:0]    io_outputs_7_payload_0_0_0_14,
  output     [7:0]    io_outputs_7_payload_0_0_0_15,
  output     [7:0]    io_outputs_7_payload_0_0_1_0,
  output     [7:0]    io_outputs_7_payload_0_0_1_1,
  output     [7:0]    io_outputs_7_payload_0_0_1_2,
  output     [7:0]    io_outputs_7_payload_0_0_1_3,
  output     [7:0]    io_outputs_7_payload_0_0_1_4,
  output     [7:0]    io_outputs_7_payload_0_0_1_5,
  output     [7:0]    io_outputs_7_payload_0_0_1_6,
  output     [7:0]    io_outputs_7_payload_0_0_1_7,
  output     [7:0]    io_outputs_7_payload_0_0_1_8,
  output     [7:0]    io_outputs_7_payload_0_0_1_9,
  output     [7:0]    io_outputs_7_payload_0_0_1_10,
  output     [7:0]    io_outputs_7_payload_0_0_1_11,
  output     [7:0]    io_outputs_7_payload_0_0_1_12,
  output     [7:0]    io_outputs_7_payload_0_0_1_13,
  output     [7:0]    io_outputs_7_payload_0_0_1_14,
  output     [7:0]    io_outputs_7_payload_0_0_1_15,
  output     [7:0]    io_outputs_7_payload_0_0_2_0,
  output     [7:0]    io_outputs_7_payload_0_0_2_1,
  output     [7:0]    io_outputs_7_payload_0_0_2_2,
  output     [7:0]    io_outputs_7_payload_0_0_2_3,
  output     [7:0]    io_outputs_7_payload_0_0_2_4,
  output     [7:0]    io_outputs_7_payload_0_0_2_5,
  output     [7:0]    io_outputs_7_payload_0_0_2_6,
  output     [7:0]    io_outputs_7_payload_0_0_2_7,
  output     [7:0]    io_outputs_7_payload_0_0_2_8,
  output     [7:0]    io_outputs_7_payload_0_0_2_9,
  output     [7:0]    io_outputs_7_payload_0_0_2_10,
  output     [7:0]    io_outputs_7_payload_0_0_2_11,
  output     [7:0]    io_outputs_7_payload_0_0_2_12,
  output     [7:0]    io_outputs_7_payload_0_0_2_13,
  output     [7:0]    io_outputs_7_payload_0_0_2_14,
  output     [7:0]    io_outputs_7_payload_0_0_2_15,
  output     [7:0]    io_outputs_7_payload_0_1_0_0,
  output     [7:0]    io_outputs_7_payload_0_1_0_1,
  output     [7:0]    io_outputs_7_payload_0_1_0_2,
  output     [7:0]    io_outputs_7_payload_0_1_0_3,
  output     [7:0]    io_outputs_7_payload_0_1_0_4,
  output     [7:0]    io_outputs_7_payload_0_1_0_5,
  output     [7:0]    io_outputs_7_payload_0_1_0_6,
  output     [7:0]    io_outputs_7_payload_0_1_0_7,
  output     [7:0]    io_outputs_7_payload_0_1_0_8,
  output     [7:0]    io_outputs_7_payload_0_1_0_9,
  output     [7:0]    io_outputs_7_payload_0_1_0_10,
  output     [7:0]    io_outputs_7_payload_0_1_0_11,
  output     [7:0]    io_outputs_7_payload_0_1_0_12,
  output     [7:0]    io_outputs_7_payload_0_1_0_13,
  output     [7:0]    io_outputs_7_payload_0_1_0_14,
  output     [7:0]    io_outputs_7_payload_0_1_0_15,
  output     [7:0]    io_outputs_7_payload_0_1_1_0,
  output     [7:0]    io_outputs_7_payload_0_1_1_1,
  output     [7:0]    io_outputs_7_payload_0_1_1_2,
  output     [7:0]    io_outputs_7_payload_0_1_1_3,
  output     [7:0]    io_outputs_7_payload_0_1_1_4,
  output     [7:0]    io_outputs_7_payload_0_1_1_5,
  output     [7:0]    io_outputs_7_payload_0_1_1_6,
  output     [7:0]    io_outputs_7_payload_0_1_1_7,
  output     [7:0]    io_outputs_7_payload_0_1_1_8,
  output     [7:0]    io_outputs_7_payload_0_1_1_9,
  output     [7:0]    io_outputs_7_payload_0_1_1_10,
  output     [7:0]    io_outputs_7_payload_0_1_1_11,
  output     [7:0]    io_outputs_7_payload_0_1_1_12,
  output     [7:0]    io_outputs_7_payload_0_1_1_13,
  output     [7:0]    io_outputs_7_payload_0_1_1_14,
  output     [7:0]    io_outputs_7_payload_0_1_1_15,
  output     [7:0]    io_outputs_7_payload_0_1_2_0,
  output     [7:0]    io_outputs_7_payload_0_1_2_1,
  output     [7:0]    io_outputs_7_payload_0_1_2_2,
  output     [7:0]    io_outputs_7_payload_0_1_2_3,
  output     [7:0]    io_outputs_7_payload_0_1_2_4,
  output     [7:0]    io_outputs_7_payload_0_1_2_5,
  output     [7:0]    io_outputs_7_payload_0_1_2_6,
  output     [7:0]    io_outputs_7_payload_0_1_2_7,
  output     [7:0]    io_outputs_7_payload_0_1_2_8,
  output     [7:0]    io_outputs_7_payload_0_1_2_9,
  output     [7:0]    io_outputs_7_payload_0_1_2_10,
  output     [7:0]    io_outputs_7_payload_0_1_2_11,
  output     [7:0]    io_outputs_7_payload_0_1_2_12,
  output     [7:0]    io_outputs_7_payload_0_1_2_13,
  output     [7:0]    io_outputs_7_payload_0_1_2_14,
  output     [7:0]    io_outputs_7_payload_0_1_2_15,
  output     [7:0]    io_outputs_7_payload_0_2_0_0,
  output     [7:0]    io_outputs_7_payload_0_2_0_1,
  output     [7:0]    io_outputs_7_payload_0_2_0_2,
  output     [7:0]    io_outputs_7_payload_0_2_0_3,
  output     [7:0]    io_outputs_7_payload_0_2_0_4,
  output     [7:0]    io_outputs_7_payload_0_2_0_5,
  output     [7:0]    io_outputs_7_payload_0_2_0_6,
  output     [7:0]    io_outputs_7_payload_0_2_0_7,
  output     [7:0]    io_outputs_7_payload_0_2_0_8,
  output     [7:0]    io_outputs_7_payload_0_2_0_9,
  output     [7:0]    io_outputs_7_payload_0_2_0_10,
  output     [7:0]    io_outputs_7_payload_0_2_0_11,
  output     [7:0]    io_outputs_7_payload_0_2_0_12,
  output     [7:0]    io_outputs_7_payload_0_2_0_13,
  output     [7:0]    io_outputs_7_payload_0_2_0_14,
  output     [7:0]    io_outputs_7_payload_0_2_0_15,
  output     [7:0]    io_outputs_7_payload_0_2_1_0,
  output     [7:0]    io_outputs_7_payload_0_2_1_1,
  output     [7:0]    io_outputs_7_payload_0_2_1_2,
  output     [7:0]    io_outputs_7_payload_0_2_1_3,
  output     [7:0]    io_outputs_7_payload_0_2_1_4,
  output     [7:0]    io_outputs_7_payload_0_2_1_5,
  output     [7:0]    io_outputs_7_payload_0_2_1_6,
  output     [7:0]    io_outputs_7_payload_0_2_1_7,
  output     [7:0]    io_outputs_7_payload_0_2_1_8,
  output     [7:0]    io_outputs_7_payload_0_2_1_9,
  output     [7:0]    io_outputs_7_payload_0_2_1_10,
  output     [7:0]    io_outputs_7_payload_0_2_1_11,
  output     [7:0]    io_outputs_7_payload_0_2_1_12,
  output     [7:0]    io_outputs_7_payload_0_2_1_13,
  output     [7:0]    io_outputs_7_payload_0_2_1_14,
  output     [7:0]    io_outputs_7_payload_0_2_1_15,
  output     [7:0]    io_outputs_7_payload_0_2_2_0,
  output     [7:0]    io_outputs_7_payload_0_2_2_1,
  output     [7:0]    io_outputs_7_payload_0_2_2_2,
  output     [7:0]    io_outputs_7_payload_0_2_2_3,
  output     [7:0]    io_outputs_7_payload_0_2_2_4,
  output     [7:0]    io_outputs_7_payload_0_2_2_5,
  output     [7:0]    io_outputs_7_payload_0_2_2_6,
  output     [7:0]    io_outputs_7_payload_0_2_2_7,
  output     [7:0]    io_outputs_7_payload_0_2_2_8,
  output     [7:0]    io_outputs_7_payload_0_2_2_9,
  output     [7:0]    io_outputs_7_payload_0_2_2_10,
  output     [7:0]    io_outputs_7_payload_0_2_2_11,
  output     [7:0]    io_outputs_7_payload_0_2_2_12,
  output     [7:0]    io_outputs_7_payload_0_2_2_13,
  output     [7:0]    io_outputs_7_payload_0_2_2_14,
  output     [7:0]    io_outputs_7_payload_0_2_2_15,
  output     [7:0]    io_outputs_7_payload_1_0_0_0,
  output     [7:0]    io_outputs_7_payload_1_0_0_1,
  output     [7:0]    io_outputs_7_payload_1_0_0_2,
  output     [7:0]    io_outputs_7_payload_1_0_0_3,
  output     [7:0]    io_outputs_7_payload_1_0_0_4,
  output     [7:0]    io_outputs_7_payload_1_0_0_5,
  output     [7:0]    io_outputs_7_payload_1_0_0_6,
  output     [7:0]    io_outputs_7_payload_1_0_0_7,
  output     [7:0]    io_outputs_7_payload_1_0_0_8,
  output     [7:0]    io_outputs_7_payload_1_0_0_9,
  output     [7:0]    io_outputs_7_payload_1_0_0_10,
  output     [7:0]    io_outputs_7_payload_1_0_0_11,
  output     [7:0]    io_outputs_7_payload_1_0_0_12,
  output     [7:0]    io_outputs_7_payload_1_0_0_13,
  output     [7:0]    io_outputs_7_payload_1_0_0_14,
  output     [7:0]    io_outputs_7_payload_1_0_0_15,
  output     [7:0]    io_outputs_7_payload_1_0_1_0,
  output     [7:0]    io_outputs_7_payload_1_0_1_1,
  output     [7:0]    io_outputs_7_payload_1_0_1_2,
  output     [7:0]    io_outputs_7_payload_1_0_1_3,
  output     [7:0]    io_outputs_7_payload_1_0_1_4,
  output     [7:0]    io_outputs_7_payload_1_0_1_5,
  output     [7:0]    io_outputs_7_payload_1_0_1_6,
  output     [7:0]    io_outputs_7_payload_1_0_1_7,
  output     [7:0]    io_outputs_7_payload_1_0_1_8,
  output     [7:0]    io_outputs_7_payload_1_0_1_9,
  output     [7:0]    io_outputs_7_payload_1_0_1_10,
  output     [7:0]    io_outputs_7_payload_1_0_1_11,
  output     [7:0]    io_outputs_7_payload_1_0_1_12,
  output     [7:0]    io_outputs_7_payload_1_0_1_13,
  output     [7:0]    io_outputs_7_payload_1_0_1_14,
  output     [7:0]    io_outputs_7_payload_1_0_1_15,
  output     [7:0]    io_outputs_7_payload_1_0_2_0,
  output     [7:0]    io_outputs_7_payload_1_0_2_1,
  output     [7:0]    io_outputs_7_payload_1_0_2_2,
  output     [7:0]    io_outputs_7_payload_1_0_2_3,
  output     [7:0]    io_outputs_7_payload_1_0_2_4,
  output     [7:0]    io_outputs_7_payload_1_0_2_5,
  output     [7:0]    io_outputs_7_payload_1_0_2_6,
  output     [7:0]    io_outputs_7_payload_1_0_2_7,
  output     [7:0]    io_outputs_7_payload_1_0_2_8,
  output     [7:0]    io_outputs_7_payload_1_0_2_9,
  output     [7:0]    io_outputs_7_payload_1_0_2_10,
  output     [7:0]    io_outputs_7_payload_1_0_2_11,
  output     [7:0]    io_outputs_7_payload_1_0_2_12,
  output     [7:0]    io_outputs_7_payload_1_0_2_13,
  output     [7:0]    io_outputs_7_payload_1_0_2_14,
  output     [7:0]    io_outputs_7_payload_1_0_2_15,
  output     [7:0]    io_outputs_7_payload_1_1_0_0,
  output     [7:0]    io_outputs_7_payload_1_1_0_1,
  output     [7:0]    io_outputs_7_payload_1_1_0_2,
  output     [7:0]    io_outputs_7_payload_1_1_0_3,
  output     [7:0]    io_outputs_7_payload_1_1_0_4,
  output     [7:0]    io_outputs_7_payload_1_1_0_5,
  output     [7:0]    io_outputs_7_payload_1_1_0_6,
  output     [7:0]    io_outputs_7_payload_1_1_0_7,
  output     [7:0]    io_outputs_7_payload_1_1_0_8,
  output     [7:0]    io_outputs_7_payload_1_1_0_9,
  output     [7:0]    io_outputs_7_payload_1_1_0_10,
  output     [7:0]    io_outputs_7_payload_1_1_0_11,
  output     [7:0]    io_outputs_7_payload_1_1_0_12,
  output     [7:0]    io_outputs_7_payload_1_1_0_13,
  output     [7:0]    io_outputs_7_payload_1_1_0_14,
  output     [7:0]    io_outputs_7_payload_1_1_0_15,
  output     [7:0]    io_outputs_7_payload_1_1_1_0,
  output     [7:0]    io_outputs_7_payload_1_1_1_1,
  output     [7:0]    io_outputs_7_payload_1_1_1_2,
  output     [7:0]    io_outputs_7_payload_1_1_1_3,
  output     [7:0]    io_outputs_7_payload_1_1_1_4,
  output     [7:0]    io_outputs_7_payload_1_1_1_5,
  output     [7:0]    io_outputs_7_payload_1_1_1_6,
  output     [7:0]    io_outputs_7_payload_1_1_1_7,
  output     [7:0]    io_outputs_7_payload_1_1_1_8,
  output     [7:0]    io_outputs_7_payload_1_1_1_9,
  output     [7:0]    io_outputs_7_payload_1_1_1_10,
  output     [7:0]    io_outputs_7_payload_1_1_1_11,
  output     [7:0]    io_outputs_7_payload_1_1_1_12,
  output     [7:0]    io_outputs_7_payload_1_1_1_13,
  output     [7:0]    io_outputs_7_payload_1_1_1_14,
  output     [7:0]    io_outputs_7_payload_1_1_1_15,
  output     [7:0]    io_outputs_7_payload_1_1_2_0,
  output     [7:0]    io_outputs_7_payload_1_1_2_1,
  output     [7:0]    io_outputs_7_payload_1_1_2_2,
  output     [7:0]    io_outputs_7_payload_1_1_2_3,
  output     [7:0]    io_outputs_7_payload_1_1_2_4,
  output     [7:0]    io_outputs_7_payload_1_1_2_5,
  output     [7:0]    io_outputs_7_payload_1_1_2_6,
  output     [7:0]    io_outputs_7_payload_1_1_2_7,
  output     [7:0]    io_outputs_7_payload_1_1_2_8,
  output     [7:0]    io_outputs_7_payload_1_1_2_9,
  output     [7:0]    io_outputs_7_payload_1_1_2_10,
  output     [7:0]    io_outputs_7_payload_1_1_2_11,
  output     [7:0]    io_outputs_7_payload_1_1_2_12,
  output     [7:0]    io_outputs_7_payload_1_1_2_13,
  output     [7:0]    io_outputs_7_payload_1_1_2_14,
  output     [7:0]    io_outputs_7_payload_1_1_2_15,
  output     [7:0]    io_outputs_7_payload_1_2_0_0,
  output     [7:0]    io_outputs_7_payload_1_2_0_1,
  output     [7:0]    io_outputs_7_payload_1_2_0_2,
  output     [7:0]    io_outputs_7_payload_1_2_0_3,
  output     [7:0]    io_outputs_7_payload_1_2_0_4,
  output     [7:0]    io_outputs_7_payload_1_2_0_5,
  output     [7:0]    io_outputs_7_payload_1_2_0_6,
  output     [7:0]    io_outputs_7_payload_1_2_0_7,
  output     [7:0]    io_outputs_7_payload_1_2_0_8,
  output     [7:0]    io_outputs_7_payload_1_2_0_9,
  output     [7:0]    io_outputs_7_payload_1_2_0_10,
  output     [7:0]    io_outputs_7_payload_1_2_0_11,
  output     [7:0]    io_outputs_7_payload_1_2_0_12,
  output     [7:0]    io_outputs_7_payload_1_2_0_13,
  output     [7:0]    io_outputs_7_payload_1_2_0_14,
  output     [7:0]    io_outputs_7_payload_1_2_0_15,
  output     [7:0]    io_outputs_7_payload_1_2_1_0,
  output     [7:0]    io_outputs_7_payload_1_2_1_1,
  output     [7:0]    io_outputs_7_payload_1_2_1_2,
  output     [7:0]    io_outputs_7_payload_1_2_1_3,
  output     [7:0]    io_outputs_7_payload_1_2_1_4,
  output     [7:0]    io_outputs_7_payload_1_2_1_5,
  output     [7:0]    io_outputs_7_payload_1_2_1_6,
  output     [7:0]    io_outputs_7_payload_1_2_1_7,
  output     [7:0]    io_outputs_7_payload_1_2_1_8,
  output     [7:0]    io_outputs_7_payload_1_2_1_9,
  output     [7:0]    io_outputs_7_payload_1_2_1_10,
  output     [7:0]    io_outputs_7_payload_1_2_1_11,
  output     [7:0]    io_outputs_7_payload_1_2_1_12,
  output     [7:0]    io_outputs_7_payload_1_2_1_13,
  output     [7:0]    io_outputs_7_payload_1_2_1_14,
  output     [7:0]    io_outputs_7_payload_1_2_1_15,
  output     [7:0]    io_outputs_7_payload_1_2_2_0,
  output     [7:0]    io_outputs_7_payload_1_2_2_1,
  output     [7:0]    io_outputs_7_payload_1_2_2_2,
  output     [7:0]    io_outputs_7_payload_1_2_2_3,
  output     [7:0]    io_outputs_7_payload_1_2_2_4,
  output     [7:0]    io_outputs_7_payload_1_2_2_5,
  output     [7:0]    io_outputs_7_payload_1_2_2_6,
  output     [7:0]    io_outputs_7_payload_1_2_2_7,
  output     [7:0]    io_outputs_7_payload_1_2_2_8,
  output     [7:0]    io_outputs_7_payload_1_2_2_9,
  output     [7:0]    io_outputs_7_payload_1_2_2_10,
  output     [7:0]    io_outputs_7_payload_1_2_2_11,
  output     [7:0]    io_outputs_7_payload_1_2_2_12,
  output     [7:0]    io_outputs_7_payload_1_2_2_13,
  output     [7:0]    io_outputs_7_payload_1_2_2_14,
  output     [7:0]    io_outputs_7_payload_1_2_2_15
);

  wire                when_Stream_l764;
  wire                when_Stream_l764_1;
  wire                when_Stream_l764_2;
  wire                when_Stream_l764_3;
  wire                when_Stream_l764_4;
  wire                when_Stream_l764_5;
  wire                when_Stream_l764_6;
  wire                when_Stream_l764_7;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l764) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l764_1) begin
      io_input_ready = io_outputs_1_ready;
    end
    if(!when_Stream_l764_2) begin
      io_input_ready = io_outputs_2_ready;
    end
    if(!when_Stream_l764_3) begin
      io_input_ready = io_outputs_3_ready;
    end
    if(!when_Stream_l764_4) begin
      io_input_ready = io_outputs_4_ready;
    end
    if(!when_Stream_l764_5) begin
      io_input_ready = io_outputs_5_ready;
    end
    if(!when_Stream_l764_6) begin
      io_input_ready = io_outputs_6_ready;
    end
    if(!when_Stream_l764_7) begin
      io_input_ready = io_outputs_7_ready;
    end
  end

  assign io_outputs_0_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_0_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_0_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_0_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_0_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_0_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_0_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_0_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_0_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_0_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_0_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_0_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_0_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_0_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_0_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_0_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_0_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_0_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_0_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_0_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_0_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_0_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_0_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_0_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_0_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_0_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_0_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_0_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_0_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_0_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_0_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_0_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_0_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_0_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_0_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_0_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_0_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_0_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_0_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_0_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_0_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_0_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_0_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_0_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_0_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_0_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_0_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_0_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_0_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_0_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_0_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_0_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_0_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_0_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_0_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_0_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_0_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_0_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_0_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_0_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_0_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_0_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_0_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_0_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_0_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_0_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_0_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_0_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_0_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_0_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_0_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_0_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_0_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_0_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_0_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_0_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_0_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_0_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_0_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_0_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_0_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_0_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_0_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_0_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_0_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_0_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_0_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_0_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_0_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_0_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_0_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_0_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_0_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_0_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_0_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_0_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_0_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_0_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_0_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_0_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_0_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_0_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_0_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_0_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_0_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_0_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_0_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_0_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_0_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_0_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_0_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_0_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_0_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_0_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_0_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_0_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_0_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_0_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_0_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_0_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_0_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_0_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_0_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_0_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_0_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_0_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_0_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_0_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_0_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_0_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_0_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_0_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_0_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_0_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_0_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_0_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_0_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_0_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_0_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_0_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_0_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_0_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_0_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_0_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_0_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_0_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_0_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_0_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_0_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_0_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_0_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_0_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_0_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_0_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_0_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_0_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_0_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_0_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_0_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_0_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_0_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_0_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_0_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_0_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_0_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_0_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_0_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_0_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_0_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_0_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_0_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_0_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_0_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_0_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_0_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_0_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_0_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_0_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_0_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_0_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_0_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_0_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_0_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_0_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_0_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_0_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_0_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_0_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_0_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_0_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_0_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_0_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_0_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_0_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_0_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_0_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_0_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_0_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_0_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_0_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_0_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_0_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_0_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_0_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_0_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_0_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_0_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_0_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_0_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_0_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_0_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_0_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_0_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_0_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_0_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_0_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_0_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_0_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_0_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_0_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_0_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_0_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_0_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_0_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_0_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_0_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_0_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_0_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_0_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_0_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_0_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_0_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_0_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_0_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_0_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_0_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_0_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_0_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_0_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_0_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_0_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_0_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_0_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_0_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_0_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_0_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_0_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_0_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_0_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_0_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_0_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_0_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_0_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_0_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_0_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_0_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_0_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_0_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_0_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_0_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_0_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_0_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_0_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_0_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_0_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_0_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_0_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_0_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_0_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_0_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_0_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_0_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_0_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_0_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_0_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_0_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_0_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_0_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_0_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_0_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_0_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_0_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_0_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_0_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_0_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_0_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_0_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_0_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764 = (3'b000 != io_select);
  always @(*) begin
    if(when_Stream_l764) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_1_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_1_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_1_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_1_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_1_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_1_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_1_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_1_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_1_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_1_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_1_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_1_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_1_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_1_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_1_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_1_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_1_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_1_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_1_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_1_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_1_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_1_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_1_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_1_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_1_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_1_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_1_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_1_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_1_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_1_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_1_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_1_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_1_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_1_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_1_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_1_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_1_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_1_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_1_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_1_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_1_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_1_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_1_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_1_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_1_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_1_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_1_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_1_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_1_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_1_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_1_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_1_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_1_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_1_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_1_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_1_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_1_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_1_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_1_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_1_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_1_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_1_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_1_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_1_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_1_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_1_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_1_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_1_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_1_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_1_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_1_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_1_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_1_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_1_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_1_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_1_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_1_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_1_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_1_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_1_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_1_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_1_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_1_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_1_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_1_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_1_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_1_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_1_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_1_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_1_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_1_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_1_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_1_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_1_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_1_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_1_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_1_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_1_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_1_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_1_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_1_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_1_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_1_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_1_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_1_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_1_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_1_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_1_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_1_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_1_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_1_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_1_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_1_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_1_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_1_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_1_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_1_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_1_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_1_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_1_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_1_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_1_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_1_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_1_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_1_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_1_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_1_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_1_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_1_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_1_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_1_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_1_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_1_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_1_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_1_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_1_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_1_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_1_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_1_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_1_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_1_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_1_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_1_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_1_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_1_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_1_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_1_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_1_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_1_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_1_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_1_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_1_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_1_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_1_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_1_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_1_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_1_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_1_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_1_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_1_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_1_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_1_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_1_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_1_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_1_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_1_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_1_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_1_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_1_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_1_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_1_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_1_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_1_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_1_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_1_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_1_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_1_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_1_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_1_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_1_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_1_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_1_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_1_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_1_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_1_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_1_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_1_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_1_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_1_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_1_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_1_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_1_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_1_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_1_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_1_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_1_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_1_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_1_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_1_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_1_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_1_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_1_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_1_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_1_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_1_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_1_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_1_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_1_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_1_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_1_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_1_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_1_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_1_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_1_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_1_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_1_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_1_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_1_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_1_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_1_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_1_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_1_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_1_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_1_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_1_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_1_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_1_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_1_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_1_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_1_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_1_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_1_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_1_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_1_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_1_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_1_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_1_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_1_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_1_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_1_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_1_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_1_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_1_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_1_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_1_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_1_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_1_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_1_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_1_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_1_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_1_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_1_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_1_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_1_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_1_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_1_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_1_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_1_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_1_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_1_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_1_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_1_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_1_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_1_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_1_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_1_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_1_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_1_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_1_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_1_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_1_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_1_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_1_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_1_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_1_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_1_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_1_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_1_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_1_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_1_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_1_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_1_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_1_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_1_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_1_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_1_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_1_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_1 = (3'b001 != io_select);
  always @(*) begin
    if(when_Stream_l764_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end

  assign io_outputs_2_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_2_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_2_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_2_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_2_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_2_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_2_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_2_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_2_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_2_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_2_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_2_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_2_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_2_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_2_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_2_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_2_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_2_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_2_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_2_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_2_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_2_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_2_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_2_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_2_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_2_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_2_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_2_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_2_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_2_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_2_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_2_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_2_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_2_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_2_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_2_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_2_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_2_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_2_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_2_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_2_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_2_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_2_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_2_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_2_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_2_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_2_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_2_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_2_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_2_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_2_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_2_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_2_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_2_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_2_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_2_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_2_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_2_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_2_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_2_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_2_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_2_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_2_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_2_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_2_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_2_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_2_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_2_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_2_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_2_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_2_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_2_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_2_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_2_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_2_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_2_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_2_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_2_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_2_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_2_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_2_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_2_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_2_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_2_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_2_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_2_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_2_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_2_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_2_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_2_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_2_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_2_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_2_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_2_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_2_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_2_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_2_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_2_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_2_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_2_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_2_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_2_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_2_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_2_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_2_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_2_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_2_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_2_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_2_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_2_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_2_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_2_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_2_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_2_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_2_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_2_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_2_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_2_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_2_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_2_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_2_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_2_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_2_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_2_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_2_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_2_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_2_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_2_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_2_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_2_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_2_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_2_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_2_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_2_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_2_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_2_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_2_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_2_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_2_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_2_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_2_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_2_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_2_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_2_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_2_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_2_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_2_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_2_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_2_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_2_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_2_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_2_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_2_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_2_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_2_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_2_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_2_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_2_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_2_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_2_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_2_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_2_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_2_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_2_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_2_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_2_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_2_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_2_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_2_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_2_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_2_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_2_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_2_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_2_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_2_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_2_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_2_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_2_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_2_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_2_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_2_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_2_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_2_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_2_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_2_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_2_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_2_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_2_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_2_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_2_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_2_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_2_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_2_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_2_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_2_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_2_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_2_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_2_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_2_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_2_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_2_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_2_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_2_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_2_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_2_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_2_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_2_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_2_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_2_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_2_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_2_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_2_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_2_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_2_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_2_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_2_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_2_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_2_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_2_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_2_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_2_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_2_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_2_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_2_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_2_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_2_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_2_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_2_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_2_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_2_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_2_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_2_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_2_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_2_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_2_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_2_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_2_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_2_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_2_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_2_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_2_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_2_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_2_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_2_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_2_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_2_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_2_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_2_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_2_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_2_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_2_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_2_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_2_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_2_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_2_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_2_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_2_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_2_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_2_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_2_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_2_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_2_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_2_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_2_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_2_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_2_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_2_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_2_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_2_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_2_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_2_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_2_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_2_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_2_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_2_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_2_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_2_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_2_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_2_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_2_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_2_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_2_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_2_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_2_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_2_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_2_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_2_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_2_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_2 = (3'b010 != io_select);
  always @(*) begin
    if(when_Stream_l764_2) begin
      io_outputs_2_valid = 1'b0;
    end else begin
      io_outputs_2_valid = io_input_valid;
    end
  end

  assign io_outputs_3_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_3_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_3_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_3_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_3_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_3_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_3_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_3_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_3_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_3_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_3_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_3_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_3_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_3_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_3_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_3_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_3_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_3_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_3_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_3_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_3_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_3_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_3_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_3_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_3_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_3_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_3_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_3_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_3_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_3_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_3_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_3_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_3_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_3_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_3_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_3_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_3_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_3_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_3_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_3_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_3_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_3_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_3_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_3_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_3_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_3_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_3_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_3_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_3_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_3_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_3_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_3_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_3_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_3_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_3_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_3_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_3_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_3_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_3_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_3_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_3_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_3_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_3_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_3_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_3_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_3_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_3_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_3_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_3_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_3_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_3_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_3_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_3_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_3_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_3_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_3_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_3_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_3_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_3_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_3_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_3_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_3_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_3_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_3_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_3_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_3_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_3_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_3_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_3_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_3_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_3_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_3_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_3_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_3_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_3_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_3_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_3_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_3_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_3_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_3_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_3_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_3_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_3_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_3_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_3_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_3_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_3_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_3_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_3_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_3_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_3_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_3_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_3_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_3_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_3_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_3_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_3_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_3_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_3_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_3_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_3_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_3_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_3_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_3_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_3_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_3_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_3_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_3_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_3_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_3_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_3_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_3_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_3_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_3_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_3_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_3_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_3_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_3_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_3_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_3_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_3_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_3_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_3_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_3_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_3_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_3_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_3_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_3_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_3_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_3_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_3_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_3_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_3_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_3_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_3_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_3_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_3_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_3_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_3_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_3_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_3_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_3_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_3_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_3_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_3_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_3_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_3_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_3_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_3_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_3_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_3_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_3_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_3_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_3_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_3_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_3_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_3_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_3_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_3_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_3_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_3_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_3_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_3_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_3_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_3_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_3_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_3_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_3_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_3_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_3_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_3_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_3_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_3_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_3_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_3_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_3_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_3_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_3_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_3_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_3_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_3_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_3_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_3_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_3_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_3_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_3_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_3_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_3_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_3_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_3_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_3_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_3_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_3_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_3_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_3_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_3_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_3_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_3_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_3_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_3_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_3_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_3_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_3_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_3_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_3_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_3_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_3_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_3_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_3_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_3_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_3_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_3_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_3_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_3_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_3_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_3_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_3_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_3_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_3_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_3_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_3_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_3_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_3_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_3_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_3_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_3_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_3_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_3_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_3_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_3_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_3_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_3_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_3_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_3_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_3_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_3_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_3_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_3_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_3_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_3_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_3_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_3_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_3_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_3_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_3_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_3_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_3_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_3_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_3_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_3_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_3_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_3_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_3_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_3_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_3_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_3_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_3_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_3_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_3_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_3_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_3_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_3_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_3_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_3_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_3_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_3_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_3_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_3_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_3 = (3'b011 != io_select);
  always @(*) begin
    if(when_Stream_l764_3) begin
      io_outputs_3_valid = 1'b0;
    end else begin
      io_outputs_3_valid = io_input_valid;
    end
  end

  assign io_outputs_4_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_4_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_4_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_4_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_4_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_4_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_4_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_4_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_4_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_4_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_4_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_4_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_4_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_4_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_4_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_4_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_4_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_4_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_4_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_4_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_4_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_4_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_4_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_4_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_4_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_4_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_4_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_4_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_4_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_4_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_4_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_4_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_4_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_4_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_4_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_4_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_4_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_4_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_4_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_4_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_4_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_4_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_4_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_4_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_4_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_4_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_4_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_4_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_4_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_4_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_4_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_4_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_4_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_4_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_4_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_4_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_4_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_4_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_4_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_4_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_4_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_4_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_4_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_4_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_4_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_4_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_4_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_4_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_4_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_4_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_4_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_4_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_4_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_4_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_4_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_4_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_4_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_4_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_4_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_4_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_4_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_4_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_4_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_4_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_4_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_4_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_4_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_4_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_4_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_4_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_4_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_4_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_4_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_4_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_4_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_4_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_4_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_4_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_4_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_4_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_4_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_4_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_4_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_4_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_4_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_4_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_4_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_4_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_4_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_4_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_4_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_4_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_4_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_4_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_4_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_4_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_4_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_4_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_4_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_4_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_4_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_4_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_4_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_4_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_4_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_4_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_4_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_4_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_4_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_4_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_4_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_4_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_4_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_4_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_4_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_4_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_4_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_4_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_4_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_4_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_4_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_4_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_4_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_4_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_4_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_4_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_4_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_4_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_4_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_4_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_4_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_4_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_4_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_4_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_4_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_4_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_4_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_4_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_4_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_4_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_4_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_4_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_4_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_4_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_4_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_4_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_4_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_4_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_4_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_4_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_4_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_4_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_4_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_4_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_4_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_4_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_4_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_4_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_4_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_4_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_4_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_4_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_4_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_4_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_4_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_4_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_4_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_4_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_4_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_4_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_4_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_4_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_4_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_4_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_4_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_4_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_4_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_4_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_4_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_4_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_4_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_4_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_4_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_4_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_4_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_4_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_4_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_4_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_4_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_4_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_4_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_4_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_4_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_4_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_4_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_4_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_4_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_4_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_4_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_4_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_4_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_4_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_4_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_4_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_4_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_4_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_4_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_4_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_4_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_4_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_4_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_4_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_4_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_4_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_4_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_4_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_4_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_4_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_4_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_4_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_4_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_4_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_4_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_4_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_4_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_4_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_4_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_4_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_4_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_4_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_4_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_4_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_4_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_4_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_4_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_4_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_4_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_4_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_4_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_4_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_4_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_4_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_4_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_4_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_4_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_4_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_4_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_4_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_4_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_4_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_4_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_4_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_4_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_4_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_4_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_4_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_4_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_4_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_4_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_4_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_4_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_4_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_4_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_4_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_4_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_4_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_4_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_4_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_4 = (3'b100 != io_select);
  always @(*) begin
    if(when_Stream_l764_4) begin
      io_outputs_4_valid = 1'b0;
    end else begin
      io_outputs_4_valid = io_input_valid;
    end
  end

  assign io_outputs_5_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_5_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_5_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_5_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_5_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_5_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_5_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_5_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_5_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_5_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_5_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_5_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_5_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_5_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_5_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_5_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_5_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_5_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_5_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_5_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_5_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_5_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_5_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_5_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_5_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_5_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_5_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_5_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_5_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_5_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_5_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_5_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_5_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_5_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_5_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_5_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_5_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_5_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_5_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_5_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_5_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_5_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_5_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_5_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_5_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_5_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_5_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_5_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_5_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_5_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_5_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_5_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_5_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_5_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_5_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_5_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_5_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_5_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_5_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_5_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_5_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_5_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_5_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_5_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_5_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_5_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_5_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_5_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_5_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_5_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_5_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_5_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_5_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_5_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_5_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_5_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_5_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_5_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_5_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_5_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_5_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_5_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_5_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_5_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_5_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_5_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_5_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_5_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_5_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_5_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_5_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_5_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_5_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_5_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_5_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_5_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_5_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_5_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_5_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_5_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_5_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_5_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_5_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_5_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_5_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_5_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_5_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_5_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_5_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_5_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_5_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_5_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_5_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_5_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_5_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_5_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_5_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_5_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_5_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_5_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_5_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_5_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_5_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_5_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_5_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_5_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_5_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_5_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_5_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_5_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_5_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_5_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_5_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_5_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_5_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_5_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_5_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_5_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_5_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_5_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_5_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_5_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_5_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_5_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_5_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_5_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_5_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_5_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_5_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_5_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_5_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_5_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_5_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_5_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_5_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_5_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_5_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_5_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_5_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_5_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_5_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_5_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_5_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_5_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_5_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_5_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_5_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_5_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_5_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_5_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_5_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_5_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_5_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_5_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_5_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_5_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_5_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_5_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_5_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_5_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_5_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_5_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_5_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_5_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_5_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_5_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_5_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_5_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_5_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_5_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_5_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_5_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_5_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_5_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_5_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_5_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_5_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_5_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_5_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_5_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_5_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_5_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_5_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_5_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_5_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_5_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_5_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_5_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_5_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_5_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_5_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_5_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_5_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_5_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_5_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_5_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_5_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_5_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_5_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_5_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_5_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_5_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_5_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_5_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_5_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_5_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_5_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_5_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_5_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_5_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_5_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_5_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_5_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_5_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_5_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_5_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_5_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_5_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_5_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_5_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_5_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_5_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_5_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_5_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_5_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_5_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_5_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_5_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_5_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_5_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_5_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_5_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_5_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_5_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_5_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_5_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_5_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_5_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_5_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_5_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_5_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_5_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_5_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_5_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_5_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_5_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_5_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_5_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_5_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_5_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_5_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_5_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_5_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_5_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_5_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_5_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_5_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_5_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_5_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_5_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_5_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_5_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_5_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_5_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_5_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_5_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_5_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_5_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_5 = (3'b101 != io_select);
  always @(*) begin
    if(when_Stream_l764_5) begin
      io_outputs_5_valid = 1'b0;
    end else begin
      io_outputs_5_valid = io_input_valid;
    end
  end

  assign io_outputs_6_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_6_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_6_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_6_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_6_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_6_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_6_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_6_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_6_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_6_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_6_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_6_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_6_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_6_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_6_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_6_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_6_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_6_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_6_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_6_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_6_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_6_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_6_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_6_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_6_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_6_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_6_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_6_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_6_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_6_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_6_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_6_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_6_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_6_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_6_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_6_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_6_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_6_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_6_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_6_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_6_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_6_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_6_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_6_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_6_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_6_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_6_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_6_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_6_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_6_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_6_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_6_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_6_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_6_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_6_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_6_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_6_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_6_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_6_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_6_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_6_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_6_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_6_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_6_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_6_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_6_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_6_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_6_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_6_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_6_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_6_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_6_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_6_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_6_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_6_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_6_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_6_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_6_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_6_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_6_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_6_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_6_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_6_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_6_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_6_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_6_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_6_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_6_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_6_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_6_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_6_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_6_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_6_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_6_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_6_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_6_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_6_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_6_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_6_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_6_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_6_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_6_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_6_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_6_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_6_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_6_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_6_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_6_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_6_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_6_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_6_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_6_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_6_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_6_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_6_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_6_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_6_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_6_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_6_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_6_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_6_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_6_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_6_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_6_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_6_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_6_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_6_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_6_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_6_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_6_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_6_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_6_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_6_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_6_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_6_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_6_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_6_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_6_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_6_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_6_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_6_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_6_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_6_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_6_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_6_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_6_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_6_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_6_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_6_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_6_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_6_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_6_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_6_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_6_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_6_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_6_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_6_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_6_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_6_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_6_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_6_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_6_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_6_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_6_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_6_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_6_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_6_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_6_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_6_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_6_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_6_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_6_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_6_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_6_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_6_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_6_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_6_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_6_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_6_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_6_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_6_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_6_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_6_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_6_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_6_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_6_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_6_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_6_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_6_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_6_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_6_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_6_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_6_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_6_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_6_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_6_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_6_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_6_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_6_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_6_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_6_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_6_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_6_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_6_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_6_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_6_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_6_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_6_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_6_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_6_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_6_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_6_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_6_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_6_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_6_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_6_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_6_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_6_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_6_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_6_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_6_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_6_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_6_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_6_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_6_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_6_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_6_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_6_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_6_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_6_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_6_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_6_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_6_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_6_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_6_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_6_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_6_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_6_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_6_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_6_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_6_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_6_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_6_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_6_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_6_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_6_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_6_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_6_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_6_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_6_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_6_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_6_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_6_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_6_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_6_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_6_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_6_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_6_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_6_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_6_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_6_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_6_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_6_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_6_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_6_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_6_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_6_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_6_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_6_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_6_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_6_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_6_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_6_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_6_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_6_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_6_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_6_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_6_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_6_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_6_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_6_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_6_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_6_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_6_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_6_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_6_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_6_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_6_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_6 = (3'b110 != io_select);
  always @(*) begin
    if(when_Stream_l764_6) begin
      io_outputs_6_valid = 1'b0;
    end else begin
      io_outputs_6_valid = io_input_valid;
    end
  end

  assign io_outputs_7_payload_0_0_0_0 = io_input_payload_0_0_0_0;
  assign io_outputs_7_payload_0_0_0_1 = io_input_payload_0_0_0_1;
  assign io_outputs_7_payload_0_0_0_2 = io_input_payload_0_0_0_2;
  assign io_outputs_7_payload_0_0_0_3 = io_input_payload_0_0_0_3;
  assign io_outputs_7_payload_0_0_0_4 = io_input_payload_0_0_0_4;
  assign io_outputs_7_payload_0_0_0_5 = io_input_payload_0_0_0_5;
  assign io_outputs_7_payload_0_0_0_6 = io_input_payload_0_0_0_6;
  assign io_outputs_7_payload_0_0_0_7 = io_input_payload_0_0_0_7;
  assign io_outputs_7_payload_0_0_0_8 = io_input_payload_0_0_0_8;
  assign io_outputs_7_payload_0_0_0_9 = io_input_payload_0_0_0_9;
  assign io_outputs_7_payload_0_0_0_10 = io_input_payload_0_0_0_10;
  assign io_outputs_7_payload_0_0_0_11 = io_input_payload_0_0_0_11;
  assign io_outputs_7_payload_0_0_0_12 = io_input_payload_0_0_0_12;
  assign io_outputs_7_payload_0_0_0_13 = io_input_payload_0_0_0_13;
  assign io_outputs_7_payload_0_0_0_14 = io_input_payload_0_0_0_14;
  assign io_outputs_7_payload_0_0_0_15 = io_input_payload_0_0_0_15;
  assign io_outputs_7_payload_0_0_1_0 = io_input_payload_0_0_1_0;
  assign io_outputs_7_payload_0_0_1_1 = io_input_payload_0_0_1_1;
  assign io_outputs_7_payload_0_0_1_2 = io_input_payload_0_0_1_2;
  assign io_outputs_7_payload_0_0_1_3 = io_input_payload_0_0_1_3;
  assign io_outputs_7_payload_0_0_1_4 = io_input_payload_0_0_1_4;
  assign io_outputs_7_payload_0_0_1_5 = io_input_payload_0_0_1_5;
  assign io_outputs_7_payload_0_0_1_6 = io_input_payload_0_0_1_6;
  assign io_outputs_7_payload_0_0_1_7 = io_input_payload_0_0_1_7;
  assign io_outputs_7_payload_0_0_1_8 = io_input_payload_0_0_1_8;
  assign io_outputs_7_payload_0_0_1_9 = io_input_payload_0_0_1_9;
  assign io_outputs_7_payload_0_0_1_10 = io_input_payload_0_0_1_10;
  assign io_outputs_7_payload_0_0_1_11 = io_input_payload_0_0_1_11;
  assign io_outputs_7_payload_0_0_1_12 = io_input_payload_0_0_1_12;
  assign io_outputs_7_payload_0_0_1_13 = io_input_payload_0_0_1_13;
  assign io_outputs_7_payload_0_0_1_14 = io_input_payload_0_0_1_14;
  assign io_outputs_7_payload_0_0_1_15 = io_input_payload_0_0_1_15;
  assign io_outputs_7_payload_0_0_2_0 = io_input_payload_0_0_2_0;
  assign io_outputs_7_payload_0_0_2_1 = io_input_payload_0_0_2_1;
  assign io_outputs_7_payload_0_0_2_2 = io_input_payload_0_0_2_2;
  assign io_outputs_7_payload_0_0_2_3 = io_input_payload_0_0_2_3;
  assign io_outputs_7_payload_0_0_2_4 = io_input_payload_0_0_2_4;
  assign io_outputs_7_payload_0_0_2_5 = io_input_payload_0_0_2_5;
  assign io_outputs_7_payload_0_0_2_6 = io_input_payload_0_0_2_6;
  assign io_outputs_7_payload_0_0_2_7 = io_input_payload_0_0_2_7;
  assign io_outputs_7_payload_0_0_2_8 = io_input_payload_0_0_2_8;
  assign io_outputs_7_payload_0_0_2_9 = io_input_payload_0_0_2_9;
  assign io_outputs_7_payload_0_0_2_10 = io_input_payload_0_0_2_10;
  assign io_outputs_7_payload_0_0_2_11 = io_input_payload_0_0_2_11;
  assign io_outputs_7_payload_0_0_2_12 = io_input_payload_0_0_2_12;
  assign io_outputs_7_payload_0_0_2_13 = io_input_payload_0_0_2_13;
  assign io_outputs_7_payload_0_0_2_14 = io_input_payload_0_0_2_14;
  assign io_outputs_7_payload_0_0_2_15 = io_input_payload_0_0_2_15;
  assign io_outputs_7_payload_0_1_0_0 = io_input_payload_0_1_0_0;
  assign io_outputs_7_payload_0_1_0_1 = io_input_payload_0_1_0_1;
  assign io_outputs_7_payload_0_1_0_2 = io_input_payload_0_1_0_2;
  assign io_outputs_7_payload_0_1_0_3 = io_input_payload_0_1_0_3;
  assign io_outputs_7_payload_0_1_0_4 = io_input_payload_0_1_0_4;
  assign io_outputs_7_payload_0_1_0_5 = io_input_payload_0_1_0_5;
  assign io_outputs_7_payload_0_1_0_6 = io_input_payload_0_1_0_6;
  assign io_outputs_7_payload_0_1_0_7 = io_input_payload_0_1_0_7;
  assign io_outputs_7_payload_0_1_0_8 = io_input_payload_0_1_0_8;
  assign io_outputs_7_payload_0_1_0_9 = io_input_payload_0_1_0_9;
  assign io_outputs_7_payload_0_1_0_10 = io_input_payload_0_1_0_10;
  assign io_outputs_7_payload_0_1_0_11 = io_input_payload_0_1_0_11;
  assign io_outputs_7_payload_0_1_0_12 = io_input_payload_0_1_0_12;
  assign io_outputs_7_payload_0_1_0_13 = io_input_payload_0_1_0_13;
  assign io_outputs_7_payload_0_1_0_14 = io_input_payload_0_1_0_14;
  assign io_outputs_7_payload_0_1_0_15 = io_input_payload_0_1_0_15;
  assign io_outputs_7_payload_0_1_1_0 = io_input_payload_0_1_1_0;
  assign io_outputs_7_payload_0_1_1_1 = io_input_payload_0_1_1_1;
  assign io_outputs_7_payload_0_1_1_2 = io_input_payload_0_1_1_2;
  assign io_outputs_7_payload_0_1_1_3 = io_input_payload_0_1_1_3;
  assign io_outputs_7_payload_0_1_1_4 = io_input_payload_0_1_1_4;
  assign io_outputs_7_payload_0_1_1_5 = io_input_payload_0_1_1_5;
  assign io_outputs_7_payload_0_1_1_6 = io_input_payload_0_1_1_6;
  assign io_outputs_7_payload_0_1_1_7 = io_input_payload_0_1_1_7;
  assign io_outputs_7_payload_0_1_1_8 = io_input_payload_0_1_1_8;
  assign io_outputs_7_payload_0_1_1_9 = io_input_payload_0_1_1_9;
  assign io_outputs_7_payload_0_1_1_10 = io_input_payload_0_1_1_10;
  assign io_outputs_7_payload_0_1_1_11 = io_input_payload_0_1_1_11;
  assign io_outputs_7_payload_0_1_1_12 = io_input_payload_0_1_1_12;
  assign io_outputs_7_payload_0_1_1_13 = io_input_payload_0_1_1_13;
  assign io_outputs_7_payload_0_1_1_14 = io_input_payload_0_1_1_14;
  assign io_outputs_7_payload_0_1_1_15 = io_input_payload_0_1_1_15;
  assign io_outputs_7_payload_0_1_2_0 = io_input_payload_0_1_2_0;
  assign io_outputs_7_payload_0_1_2_1 = io_input_payload_0_1_2_1;
  assign io_outputs_7_payload_0_1_2_2 = io_input_payload_0_1_2_2;
  assign io_outputs_7_payload_0_1_2_3 = io_input_payload_0_1_2_3;
  assign io_outputs_7_payload_0_1_2_4 = io_input_payload_0_1_2_4;
  assign io_outputs_7_payload_0_1_2_5 = io_input_payload_0_1_2_5;
  assign io_outputs_7_payload_0_1_2_6 = io_input_payload_0_1_2_6;
  assign io_outputs_7_payload_0_1_2_7 = io_input_payload_0_1_2_7;
  assign io_outputs_7_payload_0_1_2_8 = io_input_payload_0_1_2_8;
  assign io_outputs_7_payload_0_1_2_9 = io_input_payload_0_1_2_9;
  assign io_outputs_7_payload_0_1_2_10 = io_input_payload_0_1_2_10;
  assign io_outputs_7_payload_0_1_2_11 = io_input_payload_0_1_2_11;
  assign io_outputs_7_payload_0_1_2_12 = io_input_payload_0_1_2_12;
  assign io_outputs_7_payload_0_1_2_13 = io_input_payload_0_1_2_13;
  assign io_outputs_7_payload_0_1_2_14 = io_input_payload_0_1_2_14;
  assign io_outputs_7_payload_0_1_2_15 = io_input_payload_0_1_2_15;
  assign io_outputs_7_payload_0_2_0_0 = io_input_payload_0_2_0_0;
  assign io_outputs_7_payload_0_2_0_1 = io_input_payload_0_2_0_1;
  assign io_outputs_7_payload_0_2_0_2 = io_input_payload_0_2_0_2;
  assign io_outputs_7_payload_0_2_0_3 = io_input_payload_0_2_0_3;
  assign io_outputs_7_payload_0_2_0_4 = io_input_payload_0_2_0_4;
  assign io_outputs_7_payload_0_2_0_5 = io_input_payload_0_2_0_5;
  assign io_outputs_7_payload_0_2_0_6 = io_input_payload_0_2_0_6;
  assign io_outputs_7_payload_0_2_0_7 = io_input_payload_0_2_0_7;
  assign io_outputs_7_payload_0_2_0_8 = io_input_payload_0_2_0_8;
  assign io_outputs_7_payload_0_2_0_9 = io_input_payload_0_2_0_9;
  assign io_outputs_7_payload_0_2_0_10 = io_input_payload_0_2_0_10;
  assign io_outputs_7_payload_0_2_0_11 = io_input_payload_0_2_0_11;
  assign io_outputs_7_payload_0_2_0_12 = io_input_payload_0_2_0_12;
  assign io_outputs_7_payload_0_2_0_13 = io_input_payload_0_2_0_13;
  assign io_outputs_7_payload_0_2_0_14 = io_input_payload_0_2_0_14;
  assign io_outputs_7_payload_0_2_0_15 = io_input_payload_0_2_0_15;
  assign io_outputs_7_payload_0_2_1_0 = io_input_payload_0_2_1_0;
  assign io_outputs_7_payload_0_2_1_1 = io_input_payload_0_2_1_1;
  assign io_outputs_7_payload_0_2_1_2 = io_input_payload_0_2_1_2;
  assign io_outputs_7_payload_0_2_1_3 = io_input_payload_0_2_1_3;
  assign io_outputs_7_payload_0_2_1_4 = io_input_payload_0_2_1_4;
  assign io_outputs_7_payload_0_2_1_5 = io_input_payload_0_2_1_5;
  assign io_outputs_7_payload_0_2_1_6 = io_input_payload_0_2_1_6;
  assign io_outputs_7_payload_0_2_1_7 = io_input_payload_0_2_1_7;
  assign io_outputs_7_payload_0_2_1_8 = io_input_payload_0_2_1_8;
  assign io_outputs_7_payload_0_2_1_9 = io_input_payload_0_2_1_9;
  assign io_outputs_7_payload_0_2_1_10 = io_input_payload_0_2_1_10;
  assign io_outputs_7_payload_0_2_1_11 = io_input_payload_0_2_1_11;
  assign io_outputs_7_payload_0_2_1_12 = io_input_payload_0_2_1_12;
  assign io_outputs_7_payload_0_2_1_13 = io_input_payload_0_2_1_13;
  assign io_outputs_7_payload_0_2_1_14 = io_input_payload_0_2_1_14;
  assign io_outputs_7_payload_0_2_1_15 = io_input_payload_0_2_1_15;
  assign io_outputs_7_payload_0_2_2_0 = io_input_payload_0_2_2_0;
  assign io_outputs_7_payload_0_2_2_1 = io_input_payload_0_2_2_1;
  assign io_outputs_7_payload_0_2_2_2 = io_input_payload_0_2_2_2;
  assign io_outputs_7_payload_0_2_2_3 = io_input_payload_0_2_2_3;
  assign io_outputs_7_payload_0_2_2_4 = io_input_payload_0_2_2_4;
  assign io_outputs_7_payload_0_2_2_5 = io_input_payload_0_2_2_5;
  assign io_outputs_7_payload_0_2_2_6 = io_input_payload_0_2_2_6;
  assign io_outputs_7_payload_0_2_2_7 = io_input_payload_0_2_2_7;
  assign io_outputs_7_payload_0_2_2_8 = io_input_payload_0_2_2_8;
  assign io_outputs_7_payload_0_2_2_9 = io_input_payload_0_2_2_9;
  assign io_outputs_7_payload_0_2_2_10 = io_input_payload_0_2_2_10;
  assign io_outputs_7_payload_0_2_2_11 = io_input_payload_0_2_2_11;
  assign io_outputs_7_payload_0_2_2_12 = io_input_payload_0_2_2_12;
  assign io_outputs_7_payload_0_2_2_13 = io_input_payload_0_2_2_13;
  assign io_outputs_7_payload_0_2_2_14 = io_input_payload_0_2_2_14;
  assign io_outputs_7_payload_0_2_2_15 = io_input_payload_0_2_2_15;
  assign io_outputs_7_payload_1_0_0_0 = io_input_payload_1_0_0_0;
  assign io_outputs_7_payload_1_0_0_1 = io_input_payload_1_0_0_1;
  assign io_outputs_7_payload_1_0_0_2 = io_input_payload_1_0_0_2;
  assign io_outputs_7_payload_1_0_0_3 = io_input_payload_1_0_0_3;
  assign io_outputs_7_payload_1_0_0_4 = io_input_payload_1_0_0_4;
  assign io_outputs_7_payload_1_0_0_5 = io_input_payload_1_0_0_5;
  assign io_outputs_7_payload_1_0_0_6 = io_input_payload_1_0_0_6;
  assign io_outputs_7_payload_1_0_0_7 = io_input_payload_1_0_0_7;
  assign io_outputs_7_payload_1_0_0_8 = io_input_payload_1_0_0_8;
  assign io_outputs_7_payload_1_0_0_9 = io_input_payload_1_0_0_9;
  assign io_outputs_7_payload_1_0_0_10 = io_input_payload_1_0_0_10;
  assign io_outputs_7_payload_1_0_0_11 = io_input_payload_1_0_0_11;
  assign io_outputs_7_payload_1_0_0_12 = io_input_payload_1_0_0_12;
  assign io_outputs_7_payload_1_0_0_13 = io_input_payload_1_0_0_13;
  assign io_outputs_7_payload_1_0_0_14 = io_input_payload_1_0_0_14;
  assign io_outputs_7_payload_1_0_0_15 = io_input_payload_1_0_0_15;
  assign io_outputs_7_payload_1_0_1_0 = io_input_payload_1_0_1_0;
  assign io_outputs_7_payload_1_0_1_1 = io_input_payload_1_0_1_1;
  assign io_outputs_7_payload_1_0_1_2 = io_input_payload_1_0_1_2;
  assign io_outputs_7_payload_1_0_1_3 = io_input_payload_1_0_1_3;
  assign io_outputs_7_payload_1_0_1_4 = io_input_payload_1_0_1_4;
  assign io_outputs_7_payload_1_0_1_5 = io_input_payload_1_0_1_5;
  assign io_outputs_7_payload_1_0_1_6 = io_input_payload_1_0_1_6;
  assign io_outputs_7_payload_1_0_1_7 = io_input_payload_1_0_1_7;
  assign io_outputs_7_payload_1_0_1_8 = io_input_payload_1_0_1_8;
  assign io_outputs_7_payload_1_0_1_9 = io_input_payload_1_0_1_9;
  assign io_outputs_7_payload_1_0_1_10 = io_input_payload_1_0_1_10;
  assign io_outputs_7_payload_1_0_1_11 = io_input_payload_1_0_1_11;
  assign io_outputs_7_payload_1_0_1_12 = io_input_payload_1_0_1_12;
  assign io_outputs_7_payload_1_0_1_13 = io_input_payload_1_0_1_13;
  assign io_outputs_7_payload_1_0_1_14 = io_input_payload_1_0_1_14;
  assign io_outputs_7_payload_1_0_1_15 = io_input_payload_1_0_1_15;
  assign io_outputs_7_payload_1_0_2_0 = io_input_payload_1_0_2_0;
  assign io_outputs_7_payload_1_0_2_1 = io_input_payload_1_0_2_1;
  assign io_outputs_7_payload_1_0_2_2 = io_input_payload_1_0_2_2;
  assign io_outputs_7_payload_1_0_2_3 = io_input_payload_1_0_2_3;
  assign io_outputs_7_payload_1_0_2_4 = io_input_payload_1_0_2_4;
  assign io_outputs_7_payload_1_0_2_5 = io_input_payload_1_0_2_5;
  assign io_outputs_7_payload_1_0_2_6 = io_input_payload_1_0_2_6;
  assign io_outputs_7_payload_1_0_2_7 = io_input_payload_1_0_2_7;
  assign io_outputs_7_payload_1_0_2_8 = io_input_payload_1_0_2_8;
  assign io_outputs_7_payload_1_0_2_9 = io_input_payload_1_0_2_9;
  assign io_outputs_7_payload_1_0_2_10 = io_input_payload_1_0_2_10;
  assign io_outputs_7_payload_1_0_2_11 = io_input_payload_1_0_2_11;
  assign io_outputs_7_payload_1_0_2_12 = io_input_payload_1_0_2_12;
  assign io_outputs_7_payload_1_0_2_13 = io_input_payload_1_0_2_13;
  assign io_outputs_7_payload_1_0_2_14 = io_input_payload_1_0_2_14;
  assign io_outputs_7_payload_1_0_2_15 = io_input_payload_1_0_2_15;
  assign io_outputs_7_payload_1_1_0_0 = io_input_payload_1_1_0_0;
  assign io_outputs_7_payload_1_1_0_1 = io_input_payload_1_1_0_1;
  assign io_outputs_7_payload_1_1_0_2 = io_input_payload_1_1_0_2;
  assign io_outputs_7_payload_1_1_0_3 = io_input_payload_1_1_0_3;
  assign io_outputs_7_payload_1_1_0_4 = io_input_payload_1_1_0_4;
  assign io_outputs_7_payload_1_1_0_5 = io_input_payload_1_1_0_5;
  assign io_outputs_7_payload_1_1_0_6 = io_input_payload_1_1_0_6;
  assign io_outputs_7_payload_1_1_0_7 = io_input_payload_1_1_0_7;
  assign io_outputs_7_payload_1_1_0_8 = io_input_payload_1_1_0_8;
  assign io_outputs_7_payload_1_1_0_9 = io_input_payload_1_1_0_9;
  assign io_outputs_7_payload_1_1_0_10 = io_input_payload_1_1_0_10;
  assign io_outputs_7_payload_1_1_0_11 = io_input_payload_1_1_0_11;
  assign io_outputs_7_payload_1_1_0_12 = io_input_payload_1_1_0_12;
  assign io_outputs_7_payload_1_1_0_13 = io_input_payload_1_1_0_13;
  assign io_outputs_7_payload_1_1_0_14 = io_input_payload_1_1_0_14;
  assign io_outputs_7_payload_1_1_0_15 = io_input_payload_1_1_0_15;
  assign io_outputs_7_payload_1_1_1_0 = io_input_payload_1_1_1_0;
  assign io_outputs_7_payload_1_1_1_1 = io_input_payload_1_1_1_1;
  assign io_outputs_7_payload_1_1_1_2 = io_input_payload_1_1_1_2;
  assign io_outputs_7_payload_1_1_1_3 = io_input_payload_1_1_1_3;
  assign io_outputs_7_payload_1_1_1_4 = io_input_payload_1_1_1_4;
  assign io_outputs_7_payload_1_1_1_5 = io_input_payload_1_1_1_5;
  assign io_outputs_7_payload_1_1_1_6 = io_input_payload_1_1_1_6;
  assign io_outputs_7_payload_1_1_1_7 = io_input_payload_1_1_1_7;
  assign io_outputs_7_payload_1_1_1_8 = io_input_payload_1_1_1_8;
  assign io_outputs_7_payload_1_1_1_9 = io_input_payload_1_1_1_9;
  assign io_outputs_7_payload_1_1_1_10 = io_input_payload_1_1_1_10;
  assign io_outputs_7_payload_1_1_1_11 = io_input_payload_1_1_1_11;
  assign io_outputs_7_payload_1_1_1_12 = io_input_payload_1_1_1_12;
  assign io_outputs_7_payload_1_1_1_13 = io_input_payload_1_1_1_13;
  assign io_outputs_7_payload_1_1_1_14 = io_input_payload_1_1_1_14;
  assign io_outputs_7_payload_1_1_1_15 = io_input_payload_1_1_1_15;
  assign io_outputs_7_payload_1_1_2_0 = io_input_payload_1_1_2_0;
  assign io_outputs_7_payload_1_1_2_1 = io_input_payload_1_1_2_1;
  assign io_outputs_7_payload_1_1_2_2 = io_input_payload_1_1_2_2;
  assign io_outputs_7_payload_1_1_2_3 = io_input_payload_1_1_2_3;
  assign io_outputs_7_payload_1_1_2_4 = io_input_payload_1_1_2_4;
  assign io_outputs_7_payload_1_1_2_5 = io_input_payload_1_1_2_5;
  assign io_outputs_7_payload_1_1_2_6 = io_input_payload_1_1_2_6;
  assign io_outputs_7_payload_1_1_2_7 = io_input_payload_1_1_2_7;
  assign io_outputs_7_payload_1_1_2_8 = io_input_payload_1_1_2_8;
  assign io_outputs_7_payload_1_1_2_9 = io_input_payload_1_1_2_9;
  assign io_outputs_7_payload_1_1_2_10 = io_input_payload_1_1_2_10;
  assign io_outputs_7_payload_1_1_2_11 = io_input_payload_1_1_2_11;
  assign io_outputs_7_payload_1_1_2_12 = io_input_payload_1_1_2_12;
  assign io_outputs_7_payload_1_1_2_13 = io_input_payload_1_1_2_13;
  assign io_outputs_7_payload_1_1_2_14 = io_input_payload_1_1_2_14;
  assign io_outputs_7_payload_1_1_2_15 = io_input_payload_1_1_2_15;
  assign io_outputs_7_payload_1_2_0_0 = io_input_payload_1_2_0_0;
  assign io_outputs_7_payload_1_2_0_1 = io_input_payload_1_2_0_1;
  assign io_outputs_7_payload_1_2_0_2 = io_input_payload_1_2_0_2;
  assign io_outputs_7_payload_1_2_0_3 = io_input_payload_1_2_0_3;
  assign io_outputs_7_payload_1_2_0_4 = io_input_payload_1_2_0_4;
  assign io_outputs_7_payload_1_2_0_5 = io_input_payload_1_2_0_5;
  assign io_outputs_7_payload_1_2_0_6 = io_input_payload_1_2_0_6;
  assign io_outputs_7_payload_1_2_0_7 = io_input_payload_1_2_0_7;
  assign io_outputs_7_payload_1_2_0_8 = io_input_payload_1_2_0_8;
  assign io_outputs_7_payload_1_2_0_9 = io_input_payload_1_2_0_9;
  assign io_outputs_7_payload_1_2_0_10 = io_input_payload_1_2_0_10;
  assign io_outputs_7_payload_1_2_0_11 = io_input_payload_1_2_0_11;
  assign io_outputs_7_payload_1_2_0_12 = io_input_payload_1_2_0_12;
  assign io_outputs_7_payload_1_2_0_13 = io_input_payload_1_2_0_13;
  assign io_outputs_7_payload_1_2_0_14 = io_input_payload_1_2_0_14;
  assign io_outputs_7_payload_1_2_0_15 = io_input_payload_1_2_0_15;
  assign io_outputs_7_payload_1_2_1_0 = io_input_payload_1_2_1_0;
  assign io_outputs_7_payload_1_2_1_1 = io_input_payload_1_2_1_1;
  assign io_outputs_7_payload_1_2_1_2 = io_input_payload_1_2_1_2;
  assign io_outputs_7_payload_1_2_1_3 = io_input_payload_1_2_1_3;
  assign io_outputs_7_payload_1_2_1_4 = io_input_payload_1_2_1_4;
  assign io_outputs_7_payload_1_2_1_5 = io_input_payload_1_2_1_5;
  assign io_outputs_7_payload_1_2_1_6 = io_input_payload_1_2_1_6;
  assign io_outputs_7_payload_1_2_1_7 = io_input_payload_1_2_1_7;
  assign io_outputs_7_payload_1_2_1_8 = io_input_payload_1_2_1_8;
  assign io_outputs_7_payload_1_2_1_9 = io_input_payload_1_2_1_9;
  assign io_outputs_7_payload_1_2_1_10 = io_input_payload_1_2_1_10;
  assign io_outputs_7_payload_1_2_1_11 = io_input_payload_1_2_1_11;
  assign io_outputs_7_payload_1_2_1_12 = io_input_payload_1_2_1_12;
  assign io_outputs_7_payload_1_2_1_13 = io_input_payload_1_2_1_13;
  assign io_outputs_7_payload_1_2_1_14 = io_input_payload_1_2_1_14;
  assign io_outputs_7_payload_1_2_1_15 = io_input_payload_1_2_1_15;
  assign io_outputs_7_payload_1_2_2_0 = io_input_payload_1_2_2_0;
  assign io_outputs_7_payload_1_2_2_1 = io_input_payload_1_2_2_1;
  assign io_outputs_7_payload_1_2_2_2 = io_input_payload_1_2_2_2;
  assign io_outputs_7_payload_1_2_2_3 = io_input_payload_1_2_2_3;
  assign io_outputs_7_payload_1_2_2_4 = io_input_payload_1_2_2_4;
  assign io_outputs_7_payload_1_2_2_5 = io_input_payload_1_2_2_5;
  assign io_outputs_7_payload_1_2_2_6 = io_input_payload_1_2_2_6;
  assign io_outputs_7_payload_1_2_2_7 = io_input_payload_1_2_2_7;
  assign io_outputs_7_payload_1_2_2_8 = io_input_payload_1_2_2_8;
  assign io_outputs_7_payload_1_2_2_9 = io_input_payload_1_2_2_9;
  assign io_outputs_7_payload_1_2_2_10 = io_input_payload_1_2_2_10;
  assign io_outputs_7_payload_1_2_2_11 = io_input_payload_1_2_2_11;
  assign io_outputs_7_payload_1_2_2_12 = io_input_payload_1_2_2_12;
  assign io_outputs_7_payload_1_2_2_13 = io_input_payload_1_2_2_13;
  assign io_outputs_7_payload_1_2_2_14 = io_input_payload_1_2_2_14;
  assign io_outputs_7_payload_1_2_2_15 = io_input_payload_1_2_2_15;
  assign when_Stream_l764_7 = (3'b111 != io_select);
  always @(*) begin
    if(when_Stream_l764_7) begin
      io_outputs_7_valid = 1'b0;
    end else begin
      io_outputs_7_valid = io_input_valid;
    end
  end


endmodule

module LookUpTable (
  input               newTable_valid,
  output              newTable_ready,
  input      [7:0]    newTable_payload,
  input               index_valid,
  output reg          index_ready,
  input      [7:0]    index_payload_0,
  input      [7:0]    index_payload_1,
  input      [7:0]    index_payload_2,
  input      [7:0]    index_payload_3,
  input      [7:0]    index_payload_4,
  input      [7:0]    index_payload_5,
  input      [7:0]    index_payload_6,
  input      [7:0]    index_payload_7,
  input      [7:0]    index_payload_8,
  input      [7:0]    index_payload_9,
  input      [7:0]    index_payload_10,
  input      [7:0]    index_payload_11,
  input      [7:0]    index_payload_12,
  input      [7:0]    index_payload_13,
  input      [7:0]    index_payload_14,
  input      [7:0]    index_payload_15,
  output              value_valid,
  input               value_ready,
  output     [7:0]    value_payload_0,
  output     [7:0]    value_payload_1,
  output     [7:0]    value_payload_2,
  output     [7:0]    value_payload_3,
  output     [7:0]    value_payload_4,
  output     [7:0]    value_payload_5,
  output     [7:0]    value_payload_6,
  output     [7:0]    value_payload_7,
  output     [7:0]    value_payload_8,
  output     [7:0]    value_payload_9,
  output     [7:0]    value_payload_10,
  output     [7:0]    value_payload_11,
  output     [7:0]    value_payload_12,
  output     [7:0]    value_payload_13,
  output     [7:0]    value_payload_14,
  output     [7:0]    value_payload_15,
  input               clk,
  input               reset
);

  reg        [7:0]    tmp_ram_port1;
  reg        [7:0]    tmp_ram_port2;
  reg        [7:0]    tmp_ram_port3;
  reg        [7:0]    tmp_ram_port4;
  reg        [7:0]    tmp_ram_port5;
  reg        [7:0]    tmp_ram_port6;
  reg        [7:0]    tmp_ram_port7;
  reg        [7:0]    tmp_ram_port8;
  reg        [7:0]    tmp_ram_port9;
  reg        [7:0]    tmp_ram_port10;
  reg        [7:0]    tmp_ram_port11;
  reg        [7:0]    tmp_ram_port12;
  reg        [7:0]    tmp_ram_port13;
  reg        [7:0]    tmp_ram_port14;
  reg        [7:0]    tmp_ram_port15;
  reg        [7:0]    tmp_ram_port16;
  wire       [7:0]    tmp_cnt_valueNext;
  wire       [0:0]    tmp_cnt_valueNext_1;
  wire                newTable_fire;
  reg                 cnt_willIncrement;
  wire                cnt_willClear;
  reg        [7:0]    cnt_valueNext;
  reg        [7:0]    cnt_value;
  wire                cnt_willOverflowIfInc;
  wire                cnt_willOverflow;
  wire                newTable_fire_1;
  wire       [7:0]    tmp_rData_0;
  wire       [7:0]    rData_0;
  wire       [7:0]    tmp_rData_1;
  wire       [7:0]    rData_1;
  wire       [7:0]    tmp_rData_2;
  wire       [7:0]    rData_2;
  wire       [7:0]    tmp_rData_3;
  wire       [7:0]    rData_3;
  wire       [7:0]    tmp_rData_4;
  wire       [7:0]    rData_4;
  wire       [7:0]    tmp_rData_5;
  wire       [7:0]    rData_5;
  wire       [7:0]    tmp_rData_6;
  wire       [7:0]    rData_6;
  wire       [7:0]    tmp_rData_7;
  wire       [7:0]    rData_7;
  wire       [7:0]    tmp_rData_8;
  wire       [7:0]    rData_8;
  wire       [7:0]    tmp_rData_9;
  wire       [7:0]    rData_9;
  wire       [7:0]    tmp_rData_10;
  wire       [7:0]    rData_10;
  wire       [7:0]    tmp_rData_11;
  wire       [7:0]    rData_11;
  wire       [7:0]    tmp_rData_12;
  wire       [7:0]    rData_12;
  wire       [7:0]    tmp_rData_13;
  wire       [7:0]    rData_13;
  wire       [7:0]    tmp_rData_14;
  wire       [7:0]    rData_14;
  wire       [7:0]    tmp_rData_15;
  wire       [7:0]    rData_15;
  reg                 rValid;
  wire                when_LookUpTable_l25;
  (* ram_style = "distributed" *) reg [7:0] ram [0:255];

  assign tmp_cnt_valueNext_1 = cnt_willIncrement;
  assign tmp_cnt_valueNext = {7'd0, tmp_cnt_valueNext_1};
  always @(posedge clk) begin
    if(newTable_fire_1) begin
      ram[cnt_value] <= newTable_payload;
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port1 <= ram[tmp_rData_0];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port2 <= ram[tmp_rData_1];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port3 <= ram[tmp_rData_2];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port4 <= ram[tmp_rData_3];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port5 <= ram[tmp_rData_4];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port6 <= ram[tmp_rData_5];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port7 <= ram[tmp_rData_6];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port8 <= ram[tmp_rData_7];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port9 <= ram[tmp_rData_8];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port10 <= ram[tmp_rData_9];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port11 <= ram[tmp_rData_10];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port12 <= ram[tmp_rData_11];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port13 <= ram[tmp_rData_12];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port14 <= ram[tmp_rData_13];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port15 <= ram[tmp_rData_14];
    end
  end

  always @(posedge clk) begin
    if(index_ready) begin
      tmp_ram_port16 <= ram[tmp_rData_15];
    end
  end

  assign newTable_fire = (newTable_valid && newTable_ready);
  always @(*) begin
    cnt_willIncrement = 1'b0;
    if(newTable_fire) begin
      cnt_willIncrement = 1'b1;
    end
  end

  assign cnt_willClear = 1'b0;
  assign cnt_willOverflowIfInc = (cnt_value == 8'hff);
  assign cnt_willOverflow = (cnt_willOverflowIfInc && cnt_willIncrement);
  always @(*) begin
    cnt_valueNext = (cnt_value + tmp_cnt_valueNext);
    if(cnt_willClear) begin
      cnt_valueNext = 8'h0;
    end
  end

  assign newTable_fire_1 = (newTable_valid && newTable_ready);
  assign newTable_ready = 1'b1;
  assign tmp_rData_0 = index_payload_0;
  assign rData_0 = tmp_ram_port1;
  assign tmp_rData_1 = index_payload_1;
  assign rData_1 = tmp_ram_port2;
  assign tmp_rData_2 = index_payload_2;
  assign rData_2 = tmp_ram_port3;
  assign tmp_rData_3 = index_payload_3;
  assign rData_3 = tmp_ram_port4;
  assign tmp_rData_4 = index_payload_4;
  assign rData_4 = tmp_ram_port5;
  assign tmp_rData_5 = index_payload_5;
  assign rData_5 = tmp_ram_port6;
  assign tmp_rData_6 = index_payload_6;
  assign rData_6 = tmp_ram_port7;
  assign tmp_rData_7 = index_payload_7;
  assign rData_7 = tmp_ram_port8;
  assign tmp_rData_8 = index_payload_8;
  assign rData_8 = tmp_ram_port9;
  assign tmp_rData_9 = index_payload_9;
  assign rData_9 = tmp_ram_port10;
  assign tmp_rData_10 = index_payload_10;
  assign rData_10 = tmp_ram_port11;
  assign tmp_rData_11 = index_payload_11;
  assign rData_11 = tmp_ram_port12;
  assign tmp_rData_12 = index_payload_12;
  assign rData_12 = tmp_ram_port13;
  assign tmp_rData_13 = index_payload_13;
  assign rData_13 = tmp_ram_port14;
  assign tmp_rData_14 = index_payload_14;
  assign rData_14 = tmp_ram_port15;
  assign tmp_rData_15 = index_payload_15;
  assign rData_15 = tmp_ram_port16;
  always @(*) begin
    index_ready = value_ready;
    if(when_LookUpTable_l25) begin
      index_ready = 1'b1;
    end
  end

  assign when_LookUpTable_l25 = (! rValid);
  assign value_valid = rValid;
  assign value_payload_0 = rData_0;
  assign value_payload_1 = rData_1;
  assign value_payload_2 = rData_2;
  assign value_payload_3 = rData_3;
  assign value_payload_4 = rData_4;
  assign value_payload_5 = rData_5;
  assign value_payload_6 = rData_6;
  assign value_payload_7 = rData_7;
  assign value_payload_8 = rData_8;
  assign value_payload_9 = rData_9;
  assign value_payload_10 = rData_10;
  assign value_payload_11 = rData_11;
  assign value_payload_12 = rData_12;
  assign value_payload_13 = rData_13;
  assign value_payload_14 = rData_14;
  assign value_payload_15 = rData_15;
  always @(posedge clk) begin
    if(reset) begin
      cnt_value <= 8'h0;
      rValid <= 1'b0;
    end else begin
      cnt_value <= cnt_valueNext;
      if(index_ready) begin
        rValid <= index_valid;
      end
    end
  end


endmodule

module VideoPooling (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  wire                window_videoIn_ready;
  wire                window_videoOut_valid;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    window_videoOut_payload_frame_line_pixel_1_1_15;
  wire                window_videoOut_payload_frame_line_endOfLine;
  wire                window_videoOut_payload_frame_endOfFrame;
  wire                window_videoOut_payload_endOfPack;
  wire                downSample_videoIn_ready;
  wire                downSample_videoOut_valid;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_0;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_1;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_2;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_3;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_4;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_5;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_6;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_7;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_8;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_9;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_10;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_11;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_12;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_13;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_14;
  wire       [7:0]    downSample_videoOut_payload_frame_line_pixel_15;
  wire                downSample_videoOut_payload_frame_line_endOfLine;
  wire                downSample_videoOut_payload_frame_endOfFrame;
  wire                downSample_videoOut_payload_endOfPack;
  wire                merge_valid;
  reg                 merge_ready;
  wire       [7:0]    merge_payload_frame_line_pixel_0_0;
  wire       [7:0]    merge_payload_frame_line_pixel_0_1;
  wire       [7:0]    merge_payload_frame_line_pixel_0_2;
  wire       [7:0]    merge_payload_frame_line_pixel_0_3;
  wire       [7:0]    merge_payload_frame_line_pixel_0_4;
  wire       [7:0]    merge_payload_frame_line_pixel_0_5;
  wire       [7:0]    merge_payload_frame_line_pixel_0_6;
  wire       [7:0]    merge_payload_frame_line_pixel_0_7;
  wire       [7:0]    merge_payload_frame_line_pixel_0_8;
  wire       [7:0]    merge_payload_frame_line_pixel_0_9;
  wire       [7:0]    merge_payload_frame_line_pixel_0_10;
  wire       [7:0]    merge_payload_frame_line_pixel_0_11;
  wire       [7:0]    merge_payload_frame_line_pixel_0_12;
  wire       [7:0]    merge_payload_frame_line_pixel_0_13;
  wire       [7:0]    merge_payload_frame_line_pixel_0_14;
  wire       [7:0]    merge_payload_frame_line_pixel_0_15;
  wire       [7:0]    merge_payload_frame_line_pixel_1_0;
  wire       [7:0]    merge_payload_frame_line_pixel_1_1;
  wire       [7:0]    merge_payload_frame_line_pixel_1_2;
  wire       [7:0]    merge_payload_frame_line_pixel_1_3;
  wire       [7:0]    merge_payload_frame_line_pixel_1_4;
  wire       [7:0]    merge_payload_frame_line_pixel_1_5;
  wire       [7:0]    merge_payload_frame_line_pixel_1_6;
  wire       [7:0]    merge_payload_frame_line_pixel_1_7;
  wire       [7:0]    merge_payload_frame_line_pixel_1_8;
  wire       [7:0]    merge_payload_frame_line_pixel_1_9;
  wire       [7:0]    merge_payload_frame_line_pixel_1_10;
  wire       [7:0]    merge_payload_frame_line_pixel_1_11;
  wire       [7:0]    merge_payload_frame_line_pixel_1_12;
  wire       [7:0]    merge_payload_frame_line_pixel_1_13;
  wire       [7:0]    merge_payload_frame_line_pixel_1_14;
  wire       [7:0]    merge_payload_frame_line_pixel_1_15;
  wire                merge_payload_frame_line_endOfLine;
  wire                merge_payload_frame_endOfFrame;
  wire                merge_payload_endOfPack;
  wire                mergePipe_valid;
  wire                mergePipe_ready;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_0;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_1;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_2;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_3;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_4;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_5;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_6;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_7;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_8;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_9;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_10;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_11;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_12;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_13;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_14;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_0_15;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_0;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_1;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_2;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_3;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_4;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_5;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_6;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_7;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_8;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_9;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_10;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_11;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_12;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_13;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_14;
  wire       [7:0]    mergePipe_payload_frame_line_pixel_1_15;
  wire                mergePipe_payload_frame_line_endOfLine;
  wire                mergePipe_payload_frame_endOfFrame;
  wire                mergePipe_payload_endOfPack;
  reg                 merge_rValid;
  reg        [7:0]    merge_rData_frame_line_pixel_0_0;
  reg        [7:0]    merge_rData_frame_line_pixel_0_1;
  reg        [7:0]    merge_rData_frame_line_pixel_0_2;
  reg        [7:0]    merge_rData_frame_line_pixel_0_3;
  reg        [7:0]    merge_rData_frame_line_pixel_0_4;
  reg        [7:0]    merge_rData_frame_line_pixel_0_5;
  reg        [7:0]    merge_rData_frame_line_pixel_0_6;
  reg        [7:0]    merge_rData_frame_line_pixel_0_7;
  reg        [7:0]    merge_rData_frame_line_pixel_0_8;
  reg        [7:0]    merge_rData_frame_line_pixel_0_9;
  reg        [7:0]    merge_rData_frame_line_pixel_0_10;
  reg        [7:0]    merge_rData_frame_line_pixel_0_11;
  reg        [7:0]    merge_rData_frame_line_pixel_0_12;
  reg        [7:0]    merge_rData_frame_line_pixel_0_13;
  reg        [7:0]    merge_rData_frame_line_pixel_0_14;
  reg        [7:0]    merge_rData_frame_line_pixel_0_15;
  reg        [7:0]    merge_rData_frame_line_pixel_1_0;
  reg        [7:0]    merge_rData_frame_line_pixel_1_1;
  reg        [7:0]    merge_rData_frame_line_pixel_1_2;
  reg        [7:0]    merge_rData_frame_line_pixel_1_3;
  reg        [7:0]    merge_rData_frame_line_pixel_1_4;
  reg        [7:0]    merge_rData_frame_line_pixel_1_5;
  reg        [7:0]    merge_rData_frame_line_pixel_1_6;
  reg        [7:0]    merge_rData_frame_line_pixel_1_7;
  reg        [7:0]    merge_rData_frame_line_pixel_1_8;
  reg        [7:0]    merge_rData_frame_line_pixel_1_9;
  reg        [7:0]    merge_rData_frame_line_pixel_1_10;
  reg        [7:0]    merge_rData_frame_line_pixel_1_11;
  reg        [7:0]    merge_rData_frame_line_pixel_1_12;
  reg        [7:0]    merge_rData_frame_line_pixel_1_13;
  reg        [7:0]    merge_rData_frame_line_pixel_1_14;
  reg        [7:0]    merge_rData_frame_line_pixel_1_15;
  reg                 merge_rData_frame_line_endOfLine;
  reg                 merge_rData_frame_endOfFrame;
  reg                 merge_rData_endOfPack;
  wire                when_Stream_l342;
  wire                bridge_valid;
  reg                 bridge_ready;
  wire       [7:0]    bridge_payload_frame_line_pixel_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_15;
  wire                bridge_payload_frame_line_endOfLine;
  wire                bridge_payload_frame_endOfFrame;
  wire                bridge_payload_endOfPack;
  wire                bridgePipe_valid;
  wire                bridgePipe_ready;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_0;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_1;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_2;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_3;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_4;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_5;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_6;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_7;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_8;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_9;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_10;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_11;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_12;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_13;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_14;
  wire       [7:0]    bridgePipe_payload_frame_line_pixel_15;
  wire                bridgePipe_payload_frame_line_endOfLine;
  wire                bridgePipe_payload_frame_endOfFrame;
  wire                bridgePipe_payload_endOfPack;
  reg                 bridge_rValid;
  reg        [7:0]    bridge_rData_frame_line_pixel_0;
  reg        [7:0]    bridge_rData_frame_line_pixel_1;
  reg        [7:0]    bridge_rData_frame_line_pixel_2;
  reg        [7:0]    bridge_rData_frame_line_pixel_3;
  reg        [7:0]    bridge_rData_frame_line_pixel_4;
  reg        [7:0]    bridge_rData_frame_line_pixel_5;
  reg        [7:0]    bridge_rData_frame_line_pixel_6;
  reg        [7:0]    bridge_rData_frame_line_pixel_7;
  reg        [7:0]    bridge_rData_frame_line_pixel_8;
  reg        [7:0]    bridge_rData_frame_line_pixel_9;
  reg        [7:0]    bridge_rData_frame_line_pixel_10;
  reg        [7:0]    bridge_rData_frame_line_pixel_11;
  reg        [7:0]    bridge_rData_frame_line_pixel_12;
  reg        [7:0]    bridge_rData_frame_line_pixel_13;
  reg        [7:0]    bridge_rData_frame_line_pixel_14;
  reg        [7:0]    bridge_rData_frame_line_pixel_15;
  reg                 bridge_rData_frame_line_endOfLine;
  reg                 bridge_rData_frame_endOfFrame;
  reg                 bridge_rData_endOfPack;
  wire                when_Stream_l342_1;

  SlidingWindowValid window (
    .videoIn_valid                               (videoIn_valid                                         ), //i
    .videoIn_ready                               (window_videoIn_ready                                  ), //o
    .videoIn_payload_frame_line_pixel_0          (videoIn_payload_frame_line_pixel_0[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_1          (videoIn_payload_frame_line_pixel_1[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_2          (videoIn_payload_frame_line_pixel_2[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_3          (videoIn_payload_frame_line_pixel_3[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_4          (videoIn_payload_frame_line_pixel_4[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_5          (videoIn_payload_frame_line_pixel_5[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_6          (videoIn_payload_frame_line_pixel_6[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_7          (videoIn_payload_frame_line_pixel_7[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_8          (videoIn_payload_frame_line_pixel_8[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_9          (videoIn_payload_frame_line_pixel_9[7:0]               ), //i
    .videoIn_payload_frame_line_pixel_10         (videoIn_payload_frame_line_pixel_10[7:0]              ), //i
    .videoIn_payload_frame_line_pixel_11         (videoIn_payload_frame_line_pixel_11[7:0]              ), //i
    .videoIn_payload_frame_line_pixel_12         (videoIn_payload_frame_line_pixel_12[7:0]              ), //i
    .videoIn_payload_frame_line_pixel_13         (videoIn_payload_frame_line_pixel_13[7:0]              ), //i
    .videoIn_payload_frame_line_pixel_14         (videoIn_payload_frame_line_pixel_14[7:0]              ), //i
    .videoIn_payload_frame_line_pixel_15         (videoIn_payload_frame_line_pixel_15[7:0]              ), //i
    .videoIn_payload_frame_line_endOfLine        (videoIn_payload_frame_line_endOfLine                  ), //i
    .videoIn_payload_frame_endOfFrame            (videoIn_payload_frame_endOfFrame                      ), //i
    .videoIn_payload_endOfPack                   (videoIn_payload_endOfPack                             ), //i
    .videoOut_valid                              (window_videoOut_valid                                 ), //o
    .videoOut_ready                              (merge_ready                                           ), //i
    .videoOut_payload_frame_line_pixel_0_0_0     (window_videoOut_payload_frame_line_pixel_0_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_1     (window_videoOut_payload_frame_line_pixel_0_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_2     (window_videoOut_payload_frame_line_pixel_0_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_3     (window_videoOut_payload_frame_line_pixel_0_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_4     (window_videoOut_payload_frame_line_pixel_0_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_5     (window_videoOut_payload_frame_line_pixel_0_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_6     (window_videoOut_payload_frame_line_pixel_0_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_7     (window_videoOut_payload_frame_line_pixel_0_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_8     (window_videoOut_payload_frame_line_pixel_0_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_9     (window_videoOut_payload_frame_line_pixel_0_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_0_10    (window_videoOut_payload_frame_line_pixel_0_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_11    (window_videoOut_payload_frame_line_pixel_0_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_12    (window_videoOut_payload_frame_line_pixel_0_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_13    (window_videoOut_payload_frame_line_pixel_0_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_14    (window_videoOut_payload_frame_line_pixel_0_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_0_15    (window_videoOut_payload_frame_line_pixel_0_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_0     (window_videoOut_payload_frame_line_pixel_0_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_1     (window_videoOut_payload_frame_line_pixel_0_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_2     (window_videoOut_payload_frame_line_pixel_0_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_3     (window_videoOut_payload_frame_line_pixel_0_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_4     (window_videoOut_payload_frame_line_pixel_0_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_5     (window_videoOut_payload_frame_line_pixel_0_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_6     (window_videoOut_payload_frame_line_pixel_0_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_7     (window_videoOut_payload_frame_line_pixel_0_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_8     (window_videoOut_payload_frame_line_pixel_0_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_9     (window_videoOut_payload_frame_line_pixel_0_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1_10    (window_videoOut_payload_frame_line_pixel_0_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_11    (window_videoOut_payload_frame_line_pixel_0_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_12    (window_videoOut_payload_frame_line_pixel_0_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_13    (window_videoOut_payload_frame_line_pixel_0_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_14    (window_videoOut_payload_frame_line_pixel_0_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_1_15    (window_videoOut_payload_frame_line_pixel_0_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_0     (window_videoOut_payload_frame_line_pixel_1_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_1     (window_videoOut_payload_frame_line_pixel_1_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_2     (window_videoOut_payload_frame_line_pixel_1_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_3     (window_videoOut_payload_frame_line_pixel_1_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_4     (window_videoOut_payload_frame_line_pixel_1_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_5     (window_videoOut_payload_frame_line_pixel_1_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_6     (window_videoOut_payload_frame_line_pixel_1_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_7     (window_videoOut_payload_frame_line_pixel_1_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_8     (window_videoOut_payload_frame_line_pixel_1_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_9     (window_videoOut_payload_frame_line_pixel_1_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_0_10    (window_videoOut_payload_frame_line_pixel_1_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_11    (window_videoOut_payload_frame_line_pixel_1_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_12    (window_videoOut_payload_frame_line_pixel_1_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_13    (window_videoOut_payload_frame_line_pixel_1_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_14    (window_videoOut_payload_frame_line_pixel_1_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0_15    (window_videoOut_payload_frame_line_pixel_1_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_0     (window_videoOut_payload_frame_line_pixel_1_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_1     (window_videoOut_payload_frame_line_pixel_1_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_2     (window_videoOut_payload_frame_line_pixel_1_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_3     (window_videoOut_payload_frame_line_pixel_1_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_4     (window_videoOut_payload_frame_line_pixel_1_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_5     (window_videoOut_payload_frame_line_pixel_1_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_6     (window_videoOut_payload_frame_line_pixel_1_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_7     (window_videoOut_payload_frame_line_pixel_1_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_8     (window_videoOut_payload_frame_line_pixel_1_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_9     (window_videoOut_payload_frame_line_pixel_1_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1_10    (window_videoOut_payload_frame_line_pixel_1_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_11    (window_videoOut_payload_frame_line_pixel_1_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_12    (window_videoOut_payload_frame_line_pixel_1_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_13    (window_videoOut_payload_frame_line_pixel_1_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_14    (window_videoOut_payload_frame_line_pixel_1_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_1_15    (window_videoOut_payload_frame_line_pixel_1_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_endOfLine       (window_videoOut_payload_frame_line_endOfLine          ), //o
    .videoOut_payload_frame_endOfFrame           (window_videoOut_payload_frame_endOfFrame              ), //o
    .videoOut_payload_endOfPack                  (window_videoOut_payload_endOfPack                     ), //o
    .clk                                         (clk                                                   ), //i
    .reset                                       (reset                                                 )  //i
  );
  VideoDownSample downSample (
    .videoIn_valid                            (bridgePipe_valid                                      ), //i
    .videoIn_ready                            (downSample_videoIn_ready                              ), //o
    .videoIn_payload_frame_line_pixel_0       (bridgePipe_payload_frame_line_pixel_0[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_1       (bridgePipe_payload_frame_line_pixel_1[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_2       (bridgePipe_payload_frame_line_pixel_2[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_3       (bridgePipe_payload_frame_line_pixel_3[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_4       (bridgePipe_payload_frame_line_pixel_4[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_5       (bridgePipe_payload_frame_line_pixel_5[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_6       (bridgePipe_payload_frame_line_pixel_6[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_7       (bridgePipe_payload_frame_line_pixel_7[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_8       (bridgePipe_payload_frame_line_pixel_8[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_9       (bridgePipe_payload_frame_line_pixel_9[7:0]            ), //i
    .videoIn_payload_frame_line_pixel_10      (bridgePipe_payload_frame_line_pixel_10[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_11      (bridgePipe_payload_frame_line_pixel_11[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_12      (bridgePipe_payload_frame_line_pixel_12[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_13      (bridgePipe_payload_frame_line_pixel_13[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_14      (bridgePipe_payload_frame_line_pixel_14[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_15      (bridgePipe_payload_frame_line_pixel_15[7:0]           ), //i
    .videoIn_payload_frame_line_endOfLine     (bridgePipe_payload_frame_line_endOfLine               ), //i
    .videoIn_payload_frame_endOfFrame         (bridgePipe_payload_frame_endOfFrame                   ), //i
    .videoIn_payload_endOfPack                (bridgePipe_payload_endOfPack                          ), //i
    .videoOut_valid                           (downSample_videoOut_valid                             ), //o
    .videoOut_ready                           (videoOut_ready                                        ), //i
    .videoOut_payload_frame_line_pixel_0      (downSample_videoOut_payload_frame_line_pixel_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1      (downSample_videoOut_payload_frame_line_pixel_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2      (downSample_videoOut_payload_frame_line_pixel_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_3      (downSample_videoOut_payload_frame_line_pixel_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_4      (downSample_videoOut_payload_frame_line_pixel_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_5      (downSample_videoOut_payload_frame_line_pixel_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_6      (downSample_videoOut_payload_frame_line_pixel_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_7      (downSample_videoOut_payload_frame_line_pixel_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_8      (downSample_videoOut_payload_frame_line_pixel_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_9      (downSample_videoOut_payload_frame_line_pixel_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_10     (downSample_videoOut_payload_frame_line_pixel_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_11     (downSample_videoOut_payload_frame_line_pixel_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_12     (downSample_videoOut_payload_frame_line_pixel_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_13     (downSample_videoOut_payload_frame_line_pixel_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_14     (downSample_videoOut_payload_frame_line_pixel_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_15     (downSample_videoOut_payload_frame_line_pixel_15[7:0]  ), //o
    .videoOut_payload_frame_line_endOfLine    (downSample_videoOut_payload_frame_line_endOfLine      ), //o
    .videoOut_payload_frame_endOfFrame        (downSample_videoOut_payload_frame_endOfFrame          ), //o
    .videoOut_payload_endOfPack               (downSample_videoOut_payload_endOfPack                 ), //o
    .clk                                      (clk                                                   ), //i
    .reset                                    (reset                                                 )  //i
  );
  assign videoIn_ready = window_videoIn_ready;
  always @(*) begin
    merge_ready = mergePipe_ready;
    if(when_Stream_l342) begin
      merge_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mergePipe_valid);
  assign mergePipe_valid = merge_rValid;
  assign mergePipe_payload_frame_line_pixel_0_0 = merge_rData_frame_line_pixel_0_0;
  assign mergePipe_payload_frame_line_pixel_0_1 = merge_rData_frame_line_pixel_0_1;
  assign mergePipe_payload_frame_line_pixel_0_2 = merge_rData_frame_line_pixel_0_2;
  assign mergePipe_payload_frame_line_pixel_0_3 = merge_rData_frame_line_pixel_0_3;
  assign mergePipe_payload_frame_line_pixel_0_4 = merge_rData_frame_line_pixel_0_4;
  assign mergePipe_payload_frame_line_pixel_0_5 = merge_rData_frame_line_pixel_0_5;
  assign mergePipe_payload_frame_line_pixel_0_6 = merge_rData_frame_line_pixel_0_6;
  assign mergePipe_payload_frame_line_pixel_0_7 = merge_rData_frame_line_pixel_0_7;
  assign mergePipe_payload_frame_line_pixel_0_8 = merge_rData_frame_line_pixel_0_8;
  assign mergePipe_payload_frame_line_pixel_0_9 = merge_rData_frame_line_pixel_0_9;
  assign mergePipe_payload_frame_line_pixel_0_10 = merge_rData_frame_line_pixel_0_10;
  assign mergePipe_payload_frame_line_pixel_0_11 = merge_rData_frame_line_pixel_0_11;
  assign mergePipe_payload_frame_line_pixel_0_12 = merge_rData_frame_line_pixel_0_12;
  assign mergePipe_payload_frame_line_pixel_0_13 = merge_rData_frame_line_pixel_0_13;
  assign mergePipe_payload_frame_line_pixel_0_14 = merge_rData_frame_line_pixel_0_14;
  assign mergePipe_payload_frame_line_pixel_0_15 = merge_rData_frame_line_pixel_0_15;
  assign mergePipe_payload_frame_line_pixel_1_0 = merge_rData_frame_line_pixel_1_0;
  assign mergePipe_payload_frame_line_pixel_1_1 = merge_rData_frame_line_pixel_1_1;
  assign mergePipe_payload_frame_line_pixel_1_2 = merge_rData_frame_line_pixel_1_2;
  assign mergePipe_payload_frame_line_pixel_1_3 = merge_rData_frame_line_pixel_1_3;
  assign mergePipe_payload_frame_line_pixel_1_4 = merge_rData_frame_line_pixel_1_4;
  assign mergePipe_payload_frame_line_pixel_1_5 = merge_rData_frame_line_pixel_1_5;
  assign mergePipe_payload_frame_line_pixel_1_6 = merge_rData_frame_line_pixel_1_6;
  assign mergePipe_payload_frame_line_pixel_1_7 = merge_rData_frame_line_pixel_1_7;
  assign mergePipe_payload_frame_line_pixel_1_8 = merge_rData_frame_line_pixel_1_8;
  assign mergePipe_payload_frame_line_pixel_1_9 = merge_rData_frame_line_pixel_1_9;
  assign mergePipe_payload_frame_line_pixel_1_10 = merge_rData_frame_line_pixel_1_10;
  assign mergePipe_payload_frame_line_pixel_1_11 = merge_rData_frame_line_pixel_1_11;
  assign mergePipe_payload_frame_line_pixel_1_12 = merge_rData_frame_line_pixel_1_12;
  assign mergePipe_payload_frame_line_pixel_1_13 = merge_rData_frame_line_pixel_1_13;
  assign mergePipe_payload_frame_line_pixel_1_14 = merge_rData_frame_line_pixel_1_14;
  assign mergePipe_payload_frame_line_pixel_1_15 = merge_rData_frame_line_pixel_1_15;
  assign mergePipe_payload_frame_line_endOfLine = merge_rData_frame_line_endOfLine;
  assign mergePipe_payload_frame_endOfFrame = merge_rData_frame_endOfFrame;
  assign mergePipe_payload_endOfPack = merge_rData_endOfPack;
  assign merge_valid = window_videoOut_valid;
  assign merge_payload_endOfPack = window_videoOut_payload_endOfPack;
  assign merge_payload_frame_endOfFrame = window_videoOut_payload_frame_endOfFrame;
  assign merge_payload_frame_line_endOfLine = window_videoOut_payload_frame_line_endOfLine;
  assign merge_payload_frame_line_pixel_0_0 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_0) < $signed(window_videoOut_payload_frame_line_pixel_0_0_0)) ? window_videoOut_payload_frame_line_pixel_0_0_0 : window_videoOut_payload_frame_line_pixel_0_1_0);
  assign merge_payload_frame_line_pixel_0_1 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_1) < $signed(window_videoOut_payload_frame_line_pixel_0_0_1)) ? window_videoOut_payload_frame_line_pixel_0_0_1 : window_videoOut_payload_frame_line_pixel_0_1_1);
  assign merge_payload_frame_line_pixel_0_2 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_2) < $signed(window_videoOut_payload_frame_line_pixel_0_0_2)) ? window_videoOut_payload_frame_line_pixel_0_0_2 : window_videoOut_payload_frame_line_pixel_0_1_2);
  assign merge_payload_frame_line_pixel_0_3 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_3) < $signed(window_videoOut_payload_frame_line_pixel_0_0_3)) ? window_videoOut_payload_frame_line_pixel_0_0_3 : window_videoOut_payload_frame_line_pixel_0_1_3);
  assign merge_payload_frame_line_pixel_0_4 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_4) < $signed(window_videoOut_payload_frame_line_pixel_0_0_4)) ? window_videoOut_payload_frame_line_pixel_0_0_4 : window_videoOut_payload_frame_line_pixel_0_1_4);
  assign merge_payload_frame_line_pixel_0_5 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_5) < $signed(window_videoOut_payload_frame_line_pixel_0_0_5)) ? window_videoOut_payload_frame_line_pixel_0_0_5 : window_videoOut_payload_frame_line_pixel_0_1_5);
  assign merge_payload_frame_line_pixel_0_6 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_6) < $signed(window_videoOut_payload_frame_line_pixel_0_0_6)) ? window_videoOut_payload_frame_line_pixel_0_0_6 : window_videoOut_payload_frame_line_pixel_0_1_6);
  assign merge_payload_frame_line_pixel_0_7 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_7) < $signed(window_videoOut_payload_frame_line_pixel_0_0_7)) ? window_videoOut_payload_frame_line_pixel_0_0_7 : window_videoOut_payload_frame_line_pixel_0_1_7);
  assign merge_payload_frame_line_pixel_0_8 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_8) < $signed(window_videoOut_payload_frame_line_pixel_0_0_8)) ? window_videoOut_payload_frame_line_pixel_0_0_8 : window_videoOut_payload_frame_line_pixel_0_1_8);
  assign merge_payload_frame_line_pixel_0_9 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_9) < $signed(window_videoOut_payload_frame_line_pixel_0_0_9)) ? window_videoOut_payload_frame_line_pixel_0_0_9 : window_videoOut_payload_frame_line_pixel_0_1_9);
  assign merge_payload_frame_line_pixel_0_10 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_10) < $signed(window_videoOut_payload_frame_line_pixel_0_0_10)) ? window_videoOut_payload_frame_line_pixel_0_0_10 : window_videoOut_payload_frame_line_pixel_0_1_10);
  assign merge_payload_frame_line_pixel_0_11 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_11) < $signed(window_videoOut_payload_frame_line_pixel_0_0_11)) ? window_videoOut_payload_frame_line_pixel_0_0_11 : window_videoOut_payload_frame_line_pixel_0_1_11);
  assign merge_payload_frame_line_pixel_0_12 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_12) < $signed(window_videoOut_payload_frame_line_pixel_0_0_12)) ? window_videoOut_payload_frame_line_pixel_0_0_12 : window_videoOut_payload_frame_line_pixel_0_1_12);
  assign merge_payload_frame_line_pixel_0_13 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_13) < $signed(window_videoOut_payload_frame_line_pixel_0_0_13)) ? window_videoOut_payload_frame_line_pixel_0_0_13 : window_videoOut_payload_frame_line_pixel_0_1_13);
  assign merge_payload_frame_line_pixel_0_14 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_14) < $signed(window_videoOut_payload_frame_line_pixel_0_0_14)) ? window_videoOut_payload_frame_line_pixel_0_0_14 : window_videoOut_payload_frame_line_pixel_0_1_14);
  assign merge_payload_frame_line_pixel_0_15 = (($signed(window_videoOut_payload_frame_line_pixel_0_1_15) < $signed(window_videoOut_payload_frame_line_pixel_0_0_15)) ? window_videoOut_payload_frame_line_pixel_0_0_15 : window_videoOut_payload_frame_line_pixel_0_1_15);
  assign merge_payload_frame_line_pixel_1_0 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_0) < $signed(window_videoOut_payload_frame_line_pixel_1_0_0)) ? window_videoOut_payload_frame_line_pixel_1_0_0 : window_videoOut_payload_frame_line_pixel_1_1_0);
  assign merge_payload_frame_line_pixel_1_1 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_1) < $signed(window_videoOut_payload_frame_line_pixel_1_0_1)) ? window_videoOut_payload_frame_line_pixel_1_0_1 : window_videoOut_payload_frame_line_pixel_1_1_1);
  assign merge_payload_frame_line_pixel_1_2 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_2) < $signed(window_videoOut_payload_frame_line_pixel_1_0_2)) ? window_videoOut_payload_frame_line_pixel_1_0_2 : window_videoOut_payload_frame_line_pixel_1_1_2);
  assign merge_payload_frame_line_pixel_1_3 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_3) < $signed(window_videoOut_payload_frame_line_pixel_1_0_3)) ? window_videoOut_payload_frame_line_pixel_1_0_3 : window_videoOut_payload_frame_line_pixel_1_1_3);
  assign merge_payload_frame_line_pixel_1_4 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_4) < $signed(window_videoOut_payload_frame_line_pixel_1_0_4)) ? window_videoOut_payload_frame_line_pixel_1_0_4 : window_videoOut_payload_frame_line_pixel_1_1_4);
  assign merge_payload_frame_line_pixel_1_5 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_5) < $signed(window_videoOut_payload_frame_line_pixel_1_0_5)) ? window_videoOut_payload_frame_line_pixel_1_0_5 : window_videoOut_payload_frame_line_pixel_1_1_5);
  assign merge_payload_frame_line_pixel_1_6 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_6) < $signed(window_videoOut_payload_frame_line_pixel_1_0_6)) ? window_videoOut_payload_frame_line_pixel_1_0_6 : window_videoOut_payload_frame_line_pixel_1_1_6);
  assign merge_payload_frame_line_pixel_1_7 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_7) < $signed(window_videoOut_payload_frame_line_pixel_1_0_7)) ? window_videoOut_payload_frame_line_pixel_1_0_7 : window_videoOut_payload_frame_line_pixel_1_1_7);
  assign merge_payload_frame_line_pixel_1_8 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_8) < $signed(window_videoOut_payload_frame_line_pixel_1_0_8)) ? window_videoOut_payload_frame_line_pixel_1_0_8 : window_videoOut_payload_frame_line_pixel_1_1_8);
  assign merge_payload_frame_line_pixel_1_9 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_9) < $signed(window_videoOut_payload_frame_line_pixel_1_0_9)) ? window_videoOut_payload_frame_line_pixel_1_0_9 : window_videoOut_payload_frame_line_pixel_1_1_9);
  assign merge_payload_frame_line_pixel_1_10 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_10) < $signed(window_videoOut_payload_frame_line_pixel_1_0_10)) ? window_videoOut_payload_frame_line_pixel_1_0_10 : window_videoOut_payload_frame_line_pixel_1_1_10);
  assign merge_payload_frame_line_pixel_1_11 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_11) < $signed(window_videoOut_payload_frame_line_pixel_1_0_11)) ? window_videoOut_payload_frame_line_pixel_1_0_11 : window_videoOut_payload_frame_line_pixel_1_1_11);
  assign merge_payload_frame_line_pixel_1_12 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_12) < $signed(window_videoOut_payload_frame_line_pixel_1_0_12)) ? window_videoOut_payload_frame_line_pixel_1_0_12 : window_videoOut_payload_frame_line_pixel_1_1_12);
  assign merge_payload_frame_line_pixel_1_13 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_13) < $signed(window_videoOut_payload_frame_line_pixel_1_0_13)) ? window_videoOut_payload_frame_line_pixel_1_0_13 : window_videoOut_payload_frame_line_pixel_1_1_13);
  assign merge_payload_frame_line_pixel_1_14 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_14) < $signed(window_videoOut_payload_frame_line_pixel_1_0_14)) ? window_videoOut_payload_frame_line_pixel_1_0_14 : window_videoOut_payload_frame_line_pixel_1_1_14);
  assign merge_payload_frame_line_pixel_1_15 = (($signed(window_videoOut_payload_frame_line_pixel_1_1_15) < $signed(window_videoOut_payload_frame_line_pixel_1_0_15)) ? window_videoOut_payload_frame_line_pixel_1_0_15 : window_videoOut_payload_frame_line_pixel_1_1_15);
  always @(*) begin
    bridge_ready = bridgePipe_ready;
    if(when_Stream_l342_1) begin
      bridge_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! bridgePipe_valid);
  assign bridgePipe_valid = bridge_rValid;
  assign bridgePipe_payload_frame_line_pixel_0 = bridge_rData_frame_line_pixel_0;
  assign bridgePipe_payload_frame_line_pixel_1 = bridge_rData_frame_line_pixel_1;
  assign bridgePipe_payload_frame_line_pixel_2 = bridge_rData_frame_line_pixel_2;
  assign bridgePipe_payload_frame_line_pixel_3 = bridge_rData_frame_line_pixel_3;
  assign bridgePipe_payload_frame_line_pixel_4 = bridge_rData_frame_line_pixel_4;
  assign bridgePipe_payload_frame_line_pixel_5 = bridge_rData_frame_line_pixel_5;
  assign bridgePipe_payload_frame_line_pixel_6 = bridge_rData_frame_line_pixel_6;
  assign bridgePipe_payload_frame_line_pixel_7 = bridge_rData_frame_line_pixel_7;
  assign bridgePipe_payload_frame_line_pixel_8 = bridge_rData_frame_line_pixel_8;
  assign bridgePipe_payload_frame_line_pixel_9 = bridge_rData_frame_line_pixel_9;
  assign bridgePipe_payload_frame_line_pixel_10 = bridge_rData_frame_line_pixel_10;
  assign bridgePipe_payload_frame_line_pixel_11 = bridge_rData_frame_line_pixel_11;
  assign bridgePipe_payload_frame_line_pixel_12 = bridge_rData_frame_line_pixel_12;
  assign bridgePipe_payload_frame_line_pixel_13 = bridge_rData_frame_line_pixel_13;
  assign bridgePipe_payload_frame_line_pixel_14 = bridge_rData_frame_line_pixel_14;
  assign bridgePipe_payload_frame_line_pixel_15 = bridge_rData_frame_line_pixel_15;
  assign bridgePipe_payload_frame_line_endOfLine = bridge_rData_frame_line_endOfLine;
  assign bridgePipe_payload_frame_endOfFrame = bridge_rData_frame_endOfFrame;
  assign bridgePipe_payload_endOfPack = bridge_rData_endOfPack;
  assign bridge_valid = mergePipe_valid;
  assign mergePipe_ready = bridge_ready;
  assign bridge_payload_endOfPack = mergePipe_payload_endOfPack;
  assign bridge_payload_frame_endOfFrame = mergePipe_payload_frame_endOfFrame;
  assign bridge_payload_frame_line_endOfLine = mergePipe_payload_frame_line_endOfLine;
  assign bridge_payload_frame_line_pixel_0 = (($signed(mergePipe_payload_frame_line_pixel_1_0) < $signed(mergePipe_payload_frame_line_pixel_0_0)) ? mergePipe_payload_frame_line_pixel_0_0 : mergePipe_payload_frame_line_pixel_1_0);
  assign bridge_payload_frame_line_pixel_1 = (($signed(mergePipe_payload_frame_line_pixel_1_1) < $signed(mergePipe_payload_frame_line_pixel_0_1)) ? mergePipe_payload_frame_line_pixel_0_1 : mergePipe_payload_frame_line_pixel_1_1);
  assign bridge_payload_frame_line_pixel_2 = (($signed(mergePipe_payload_frame_line_pixel_1_2) < $signed(mergePipe_payload_frame_line_pixel_0_2)) ? mergePipe_payload_frame_line_pixel_0_2 : mergePipe_payload_frame_line_pixel_1_2);
  assign bridge_payload_frame_line_pixel_3 = (($signed(mergePipe_payload_frame_line_pixel_1_3) < $signed(mergePipe_payload_frame_line_pixel_0_3)) ? mergePipe_payload_frame_line_pixel_0_3 : mergePipe_payload_frame_line_pixel_1_3);
  assign bridge_payload_frame_line_pixel_4 = (($signed(mergePipe_payload_frame_line_pixel_1_4) < $signed(mergePipe_payload_frame_line_pixel_0_4)) ? mergePipe_payload_frame_line_pixel_0_4 : mergePipe_payload_frame_line_pixel_1_4);
  assign bridge_payload_frame_line_pixel_5 = (($signed(mergePipe_payload_frame_line_pixel_1_5) < $signed(mergePipe_payload_frame_line_pixel_0_5)) ? mergePipe_payload_frame_line_pixel_0_5 : mergePipe_payload_frame_line_pixel_1_5);
  assign bridge_payload_frame_line_pixel_6 = (($signed(mergePipe_payload_frame_line_pixel_1_6) < $signed(mergePipe_payload_frame_line_pixel_0_6)) ? mergePipe_payload_frame_line_pixel_0_6 : mergePipe_payload_frame_line_pixel_1_6);
  assign bridge_payload_frame_line_pixel_7 = (($signed(mergePipe_payload_frame_line_pixel_1_7) < $signed(mergePipe_payload_frame_line_pixel_0_7)) ? mergePipe_payload_frame_line_pixel_0_7 : mergePipe_payload_frame_line_pixel_1_7);
  assign bridge_payload_frame_line_pixel_8 = (($signed(mergePipe_payload_frame_line_pixel_1_8) < $signed(mergePipe_payload_frame_line_pixel_0_8)) ? mergePipe_payload_frame_line_pixel_0_8 : mergePipe_payload_frame_line_pixel_1_8);
  assign bridge_payload_frame_line_pixel_9 = (($signed(mergePipe_payload_frame_line_pixel_1_9) < $signed(mergePipe_payload_frame_line_pixel_0_9)) ? mergePipe_payload_frame_line_pixel_0_9 : mergePipe_payload_frame_line_pixel_1_9);
  assign bridge_payload_frame_line_pixel_10 = (($signed(mergePipe_payload_frame_line_pixel_1_10) < $signed(mergePipe_payload_frame_line_pixel_0_10)) ? mergePipe_payload_frame_line_pixel_0_10 : mergePipe_payload_frame_line_pixel_1_10);
  assign bridge_payload_frame_line_pixel_11 = (($signed(mergePipe_payload_frame_line_pixel_1_11) < $signed(mergePipe_payload_frame_line_pixel_0_11)) ? mergePipe_payload_frame_line_pixel_0_11 : mergePipe_payload_frame_line_pixel_1_11);
  assign bridge_payload_frame_line_pixel_12 = (($signed(mergePipe_payload_frame_line_pixel_1_12) < $signed(mergePipe_payload_frame_line_pixel_0_12)) ? mergePipe_payload_frame_line_pixel_0_12 : mergePipe_payload_frame_line_pixel_1_12);
  assign bridge_payload_frame_line_pixel_13 = (($signed(mergePipe_payload_frame_line_pixel_1_13) < $signed(mergePipe_payload_frame_line_pixel_0_13)) ? mergePipe_payload_frame_line_pixel_0_13 : mergePipe_payload_frame_line_pixel_1_13);
  assign bridge_payload_frame_line_pixel_14 = (($signed(mergePipe_payload_frame_line_pixel_1_14) < $signed(mergePipe_payload_frame_line_pixel_0_14)) ? mergePipe_payload_frame_line_pixel_0_14 : mergePipe_payload_frame_line_pixel_1_14);
  assign bridge_payload_frame_line_pixel_15 = (($signed(mergePipe_payload_frame_line_pixel_1_15) < $signed(mergePipe_payload_frame_line_pixel_0_15)) ? mergePipe_payload_frame_line_pixel_0_15 : mergePipe_payload_frame_line_pixel_1_15);
  assign bridgePipe_ready = downSample_videoIn_ready;
  assign videoOut_valid = downSample_videoOut_valid;
  assign videoOut_payload_frame_line_pixel_0 = downSample_videoOut_payload_frame_line_pixel_0;
  assign videoOut_payload_frame_line_pixel_1 = downSample_videoOut_payload_frame_line_pixel_1;
  assign videoOut_payload_frame_line_pixel_2 = downSample_videoOut_payload_frame_line_pixel_2;
  assign videoOut_payload_frame_line_pixel_3 = downSample_videoOut_payload_frame_line_pixel_3;
  assign videoOut_payload_frame_line_pixel_4 = downSample_videoOut_payload_frame_line_pixel_4;
  assign videoOut_payload_frame_line_pixel_5 = downSample_videoOut_payload_frame_line_pixel_5;
  assign videoOut_payload_frame_line_pixel_6 = downSample_videoOut_payload_frame_line_pixel_6;
  assign videoOut_payload_frame_line_pixel_7 = downSample_videoOut_payload_frame_line_pixel_7;
  assign videoOut_payload_frame_line_pixel_8 = downSample_videoOut_payload_frame_line_pixel_8;
  assign videoOut_payload_frame_line_pixel_9 = downSample_videoOut_payload_frame_line_pixel_9;
  assign videoOut_payload_frame_line_pixel_10 = downSample_videoOut_payload_frame_line_pixel_10;
  assign videoOut_payload_frame_line_pixel_11 = downSample_videoOut_payload_frame_line_pixel_11;
  assign videoOut_payload_frame_line_pixel_12 = downSample_videoOut_payload_frame_line_pixel_12;
  assign videoOut_payload_frame_line_pixel_13 = downSample_videoOut_payload_frame_line_pixel_13;
  assign videoOut_payload_frame_line_pixel_14 = downSample_videoOut_payload_frame_line_pixel_14;
  assign videoOut_payload_frame_line_pixel_15 = downSample_videoOut_payload_frame_line_pixel_15;
  assign videoOut_payload_frame_line_endOfLine = downSample_videoOut_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_endOfFrame = downSample_videoOut_payload_frame_endOfFrame;
  assign videoOut_payload_endOfPack = downSample_videoOut_payload_endOfPack;
  always @(posedge clk) begin
    if(reset) begin
      merge_rValid <= 1'b0;
      bridge_rValid <= 1'b0;
    end else begin
      if(merge_ready) begin
        merge_rValid <= merge_valid;
      end
      if(bridge_ready) begin
        bridge_rValid <= bridge_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(merge_ready) begin
      merge_rData_frame_line_pixel_0_0 <= merge_payload_frame_line_pixel_0_0;
      merge_rData_frame_line_pixel_0_1 <= merge_payload_frame_line_pixel_0_1;
      merge_rData_frame_line_pixel_0_2 <= merge_payload_frame_line_pixel_0_2;
      merge_rData_frame_line_pixel_0_3 <= merge_payload_frame_line_pixel_0_3;
      merge_rData_frame_line_pixel_0_4 <= merge_payload_frame_line_pixel_0_4;
      merge_rData_frame_line_pixel_0_5 <= merge_payload_frame_line_pixel_0_5;
      merge_rData_frame_line_pixel_0_6 <= merge_payload_frame_line_pixel_0_6;
      merge_rData_frame_line_pixel_0_7 <= merge_payload_frame_line_pixel_0_7;
      merge_rData_frame_line_pixel_0_8 <= merge_payload_frame_line_pixel_0_8;
      merge_rData_frame_line_pixel_0_9 <= merge_payload_frame_line_pixel_0_9;
      merge_rData_frame_line_pixel_0_10 <= merge_payload_frame_line_pixel_0_10;
      merge_rData_frame_line_pixel_0_11 <= merge_payload_frame_line_pixel_0_11;
      merge_rData_frame_line_pixel_0_12 <= merge_payload_frame_line_pixel_0_12;
      merge_rData_frame_line_pixel_0_13 <= merge_payload_frame_line_pixel_0_13;
      merge_rData_frame_line_pixel_0_14 <= merge_payload_frame_line_pixel_0_14;
      merge_rData_frame_line_pixel_0_15 <= merge_payload_frame_line_pixel_0_15;
      merge_rData_frame_line_pixel_1_0 <= merge_payload_frame_line_pixel_1_0;
      merge_rData_frame_line_pixel_1_1 <= merge_payload_frame_line_pixel_1_1;
      merge_rData_frame_line_pixel_1_2 <= merge_payload_frame_line_pixel_1_2;
      merge_rData_frame_line_pixel_1_3 <= merge_payload_frame_line_pixel_1_3;
      merge_rData_frame_line_pixel_1_4 <= merge_payload_frame_line_pixel_1_4;
      merge_rData_frame_line_pixel_1_5 <= merge_payload_frame_line_pixel_1_5;
      merge_rData_frame_line_pixel_1_6 <= merge_payload_frame_line_pixel_1_6;
      merge_rData_frame_line_pixel_1_7 <= merge_payload_frame_line_pixel_1_7;
      merge_rData_frame_line_pixel_1_8 <= merge_payload_frame_line_pixel_1_8;
      merge_rData_frame_line_pixel_1_9 <= merge_payload_frame_line_pixel_1_9;
      merge_rData_frame_line_pixel_1_10 <= merge_payload_frame_line_pixel_1_10;
      merge_rData_frame_line_pixel_1_11 <= merge_payload_frame_line_pixel_1_11;
      merge_rData_frame_line_pixel_1_12 <= merge_payload_frame_line_pixel_1_12;
      merge_rData_frame_line_pixel_1_13 <= merge_payload_frame_line_pixel_1_13;
      merge_rData_frame_line_pixel_1_14 <= merge_payload_frame_line_pixel_1_14;
      merge_rData_frame_line_pixel_1_15 <= merge_payload_frame_line_pixel_1_15;
      merge_rData_frame_line_endOfLine <= merge_payload_frame_line_endOfLine;
      merge_rData_frame_endOfFrame <= merge_payload_frame_endOfFrame;
      merge_rData_endOfPack <= merge_payload_endOfPack;
    end
    if(bridge_ready) begin
      bridge_rData_frame_line_pixel_0 <= bridge_payload_frame_line_pixel_0;
      bridge_rData_frame_line_pixel_1 <= bridge_payload_frame_line_pixel_1;
      bridge_rData_frame_line_pixel_2 <= bridge_payload_frame_line_pixel_2;
      bridge_rData_frame_line_pixel_3 <= bridge_payload_frame_line_pixel_3;
      bridge_rData_frame_line_pixel_4 <= bridge_payload_frame_line_pixel_4;
      bridge_rData_frame_line_pixel_5 <= bridge_payload_frame_line_pixel_5;
      bridge_rData_frame_line_pixel_6 <= bridge_payload_frame_line_pixel_6;
      bridge_rData_frame_line_pixel_7 <= bridge_payload_frame_line_pixel_7;
      bridge_rData_frame_line_pixel_8 <= bridge_payload_frame_line_pixel_8;
      bridge_rData_frame_line_pixel_9 <= bridge_payload_frame_line_pixel_9;
      bridge_rData_frame_line_pixel_10 <= bridge_payload_frame_line_pixel_10;
      bridge_rData_frame_line_pixel_11 <= bridge_payload_frame_line_pixel_11;
      bridge_rData_frame_line_pixel_12 <= bridge_payload_frame_line_pixel_12;
      bridge_rData_frame_line_pixel_13 <= bridge_payload_frame_line_pixel_13;
      bridge_rData_frame_line_pixel_14 <= bridge_payload_frame_line_pixel_14;
      bridge_rData_frame_line_pixel_15 <= bridge_payload_frame_line_pixel_15;
      bridge_rData_frame_line_endOfLine <= bridge_payload_frame_line_endOfLine;
      bridge_rData_frame_endOfFrame <= bridge_payload_frame_endOfFrame;
      bridge_rData_endOfPack <= bridge_payload_endOfPack;
    end
  end


endmodule

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

//PecaUnit replaced by PecaUnit

module PecaUnit (
  input      [7:0]    numberOfInputFrames,
  input      [7:0]    numberOfOutputFrames,
  input               inputs_valid,
  output              inputs_ready,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_0,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_1,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_2,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_3,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_4,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_5,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_6,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_7,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_8,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_9,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_10,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_11,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_12,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_13,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_14,
  input      [7:0]    inputs_payload_frame_line_pixel_0_0_15,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_0,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_1,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_2,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_3,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_4,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_5,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_6,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_7,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_8,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_9,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_10,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_11,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_12,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_13,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_14,
  input      [7:0]    inputs_payload_frame_line_pixel_0_1_15,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_0,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_1,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_2,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_3,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_4,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_5,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_6,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_7,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_8,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_9,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_10,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_11,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_12,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_13,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_14,
  input      [7:0]    inputs_payload_frame_line_pixel_0_2_15,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_0,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_1,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_2,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_3,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_4,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_5,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_6,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_7,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_8,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_9,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_10,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_11,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_12,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_13,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_14,
  input      [7:0]    inputs_payload_frame_line_pixel_1_0_15,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_0,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_1,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_2,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_3,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_4,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_5,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_6,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_7,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_8,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_9,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_10,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_11,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_12,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_13,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_14,
  input      [7:0]    inputs_payload_frame_line_pixel_1_1_15,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_0,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_1,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_2,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_3,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_4,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_5,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_6,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_7,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_8,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_9,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_10,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_11,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_12,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_13,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_14,
  input      [7:0]    inputs_payload_frame_line_pixel_1_2_15,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_0,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_1,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_2,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_3,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_4,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_5,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_6,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_7,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_8,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_9,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_10,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_11,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_12,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_13,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_14,
  input      [7:0]    inputs_payload_frame_line_pixel_2_0_15,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_0,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_1,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_2,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_3,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_4,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_5,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_6,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_7,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_8,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_9,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_10,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_11,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_12,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_13,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_14,
  input      [7:0]    inputs_payload_frame_line_pixel_2_1_15,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_0,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_1,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_2,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_3,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_4,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_5,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_6,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_7,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_8,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_9,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_10,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_11,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_12,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_13,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_14,
  input      [7:0]    inputs_payload_frame_line_pixel_2_2_15,
  input               inputs_payload_frame_line_endOfLine,
  input               inputs_payload_frame_endOfFrame,
  input               inputs_payload_endOfPack,
  input               weights_valid,
  output              weights_ready,
  input      [7:0]    weights_payload_0_0_0_0,
  input      [7:0]    weights_payload_0_0_0_1,
  input      [7:0]    weights_payload_0_0_0_2,
  input      [7:0]    weights_payload_0_0_0_3,
  input      [7:0]    weights_payload_0_0_0_4,
  input      [7:0]    weights_payload_0_0_0_5,
  input      [7:0]    weights_payload_0_0_0_6,
  input      [7:0]    weights_payload_0_0_0_7,
  input      [7:0]    weights_payload_0_0_0_8,
  input      [7:0]    weights_payload_0_0_0_9,
  input      [7:0]    weights_payload_0_0_0_10,
  input      [7:0]    weights_payload_0_0_0_11,
  input      [7:0]    weights_payload_0_0_0_12,
  input      [7:0]    weights_payload_0_0_0_13,
  input      [7:0]    weights_payload_0_0_0_14,
  input      [7:0]    weights_payload_0_0_0_15,
  input      [7:0]    weights_payload_0_0_1_0,
  input      [7:0]    weights_payload_0_0_1_1,
  input      [7:0]    weights_payload_0_0_1_2,
  input      [7:0]    weights_payload_0_0_1_3,
  input      [7:0]    weights_payload_0_0_1_4,
  input      [7:0]    weights_payload_0_0_1_5,
  input      [7:0]    weights_payload_0_0_1_6,
  input      [7:0]    weights_payload_0_0_1_7,
  input      [7:0]    weights_payload_0_0_1_8,
  input      [7:0]    weights_payload_0_0_1_9,
  input      [7:0]    weights_payload_0_0_1_10,
  input      [7:0]    weights_payload_0_0_1_11,
  input      [7:0]    weights_payload_0_0_1_12,
  input      [7:0]    weights_payload_0_0_1_13,
  input      [7:0]    weights_payload_0_0_1_14,
  input      [7:0]    weights_payload_0_0_1_15,
  input      [7:0]    weights_payload_0_0_2_0,
  input      [7:0]    weights_payload_0_0_2_1,
  input      [7:0]    weights_payload_0_0_2_2,
  input      [7:0]    weights_payload_0_0_2_3,
  input      [7:0]    weights_payload_0_0_2_4,
  input      [7:0]    weights_payload_0_0_2_5,
  input      [7:0]    weights_payload_0_0_2_6,
  input      [7:0]    weights_payload_0_0_2_7,
  input      [7:0]    weights_payload_0_0_2_8,
  input      [7:0]    weights_payload_0_0_2_9,
  input      [7:0]    weights_payload_0_0_2_10,
  input      [7:0]    weights_payload_0_0_2_11,
  input      [7:0]    weights_payload_0_0_2_12,
  input      [7:0]    weights_payload_0_0_2_13,
  input      [7:0]    weights_payload_0_0_2_14,
  input      [7:0]    weights_payload_0_0_2_15,
  input      [7:0]    weights_payload_0_1_0_0,
  input      [7:0]    weights_payload_0_1_0_1,
  input      [7:0]    weights_payload_0_1_0_2,
  input      [7:0]    weights_payload_0_1_0_3,
  input      [7:0]    weights_payload_0_1_0_4,
  input      [7:0]    weights_payload_0_1_0_5,
  input      [7:0]    weights_payload_0_1_0_6,
  input      [7:0]    weights_payload_0_1_0_7,
  input      [7:0]    weights_payload_0_1_0_8,
  input      [7:0]    weights_payload_0_1_0_9,
  input      [7:0]    weights_payload_0_1_0_10,
  input      [7:0]    weights_payload_0_1_0_11,
  input      [7:0]    weights_payload_0_1_0_12,
  input      [7:0]    weights_payload_0_1_0_13,
  input      [7:0]    weights_payload_0_1_0_14,
  input      [7:0]    weights_payload_0_1_0_15,
  input      [7:0]    weights_payload_0_1_1_0,
  input      [7:0]    weights_payload_0_1_1_1,
  input      [7:0]    weights_payload_0_1_1_2,
  input      [7:0]    weights_payload_0_1_1_3,
  input      [7:0]    weights_payload_0_1_1_4,
  input      [7:0]    weights_payload_0_1_1_5,
  input      [7:0]    weights_payload_0_1_1_6,
  input      [7:0]    weights_payload_0_1_1_7,
  input      [7:0]    weights_payload_0_1_1_8,
  input      [7:0]    weights_payload_0_1_1_9,
  input      [7:0]    weights_payload_0_1_1_10,
  input      [7:0]    weights_payload_0_1_1_11,
  input      [7:0]    weights_payload_0_1_1_12,
  input      [7:0]    weights_payload_0_1_1_13,
  input      [7:0]    weights_payload_0_1_1_14,
  input      [7:0]    weights_payload_0_1_1_15,
  input      [7:0]    weights_payload_0_1_2_0,
  input      [7:0]    weights_payload_0_1_2_1,
  input      [7:0]    weights_payload_0_1_2_2,
  input      [7:0]    weights_payload_0_1_2_3,
  input      [7:0]    weights_payload_0_1_2_4,
  input      [7:0]    weights_payload_0_1_2_5,
  input      [7:0]    weights_payload_0_1_2_6,
  input      [7:0]    weights_payload_0_1_2_7,
  input      [7:0]    weights_payload_0_1_2_8,
  input      [7:0]    weights_payload_0_1_2_9,
  input      [7:0]    weights_payload_0_1_2_10,
  input      [7:0]    weights_payload_0_1_2_11,
  input      [7:0]    weights_payload_0_1_2_12,
  input      [7:0]    weights_payload_0_1_2_13,
  input      [7:0]    weights_payload_0_1_2_14,
  input      [7:0]    weights_payload_0_1_2_15,
  input      [7:0]    weights_payload_0_2_0_0,
  input      [7:0]    weights_payload_0_2_0_1,
  input      [7:0]    weights_payload_0_2_0_2,
  input      [7:0]    weights_payload_0_2_0_3,
  input      [7:0]    weights_payload_0_2_0_4,
  input      [7:0]    weights_payload_0_2_0_5,
  input      [7:0]    weights_payload_0_2_0_6,
  input      [7:0]    weights_payload_0_2_0_7,
  input      [7:0]    weights_payload_0_2_0_8,
  input      [7:0]    weights_payload_0_2_0_9,
  input      [7:0]    weights_payload_0_2_0_10,
  input      [7:0]    weights_payload_0_2_0_11,
  input      [7:0]    weights_payload_0_2_0_12,
  input      [7:0]    weights_payload_0_2_0_13,
  input      [7:0]    weights_payload_0_2_0_14,
  input      [7:0]    weights_payload_0_2_0_15,
  input      [7:0]    weights_payload_0_2_1_0,
  input      [7:0]    weights_payload_0_2_1_1,
  input      [7:0]    weights_payload_0_2_1_2,
  input      [7:0]    weights_payload_0_2_1_3,
  input      [7:0]    weights_payload_0_2_1_4,
  input      [7:0]    weights_payload_0_2_1_5,
  input      [7:0]    weights_payload_0_2_1_6,
  input      [7:0]    weights_payload_0_2_1_7,
  input      [7:0]    weights_payload_0_2_1_8,
  input      [7:0]    weights_payload_0_2_1_9,
  input      [7:0]    weights_payload_0_2_1_10,
  input      [7:0]    weights_payload_0_2_1_11,
  input      [7:0]    weights_payload_0_2_1_12,
  input      [7:0]    weights_payload_0_2_1_13,
  input      [7:0]    weights_payload_0_2_1_14,
  input      [7:0]    weights_payload_0_2_1_15,
  input      [7:0]    weights_payload_0_2_2_0,
  input      [7:0]    weights_payload_0_2_2_1,
  input      [7:0]    weights_payload_0_2_2_2,
  input      [7:0]    weights_payload_0_2_2_3,
  input      [7:0]    weights_payload_0_2_2_4,
  input      [7:0]    weights_payload_0_2_2_5,
  input      [7:0]    weights_payload_0_2_2_6,
  input      [7:0]    weights_payload_0_2_2_7,
  input      [7:0]    weights_payload_0_2_2_8,
  input      [7:0]    weights_payload_0_2_2_9,
  input      [7:0]    weights_payload_0_2_2_10,
  input      [7:0]    weights_payload_0_2_2_11,
  input      [7:0]    weights_payload_0_2_2_12,
  input      [7:0]    weights_payload_0_2_2_13,
  input      [7:0]    weights_payload_0_2_2_14,
  input      [7:0]    weights_payload_0_2_2_15,
  input      [7:0]    weights_payload_1_0_0_0,
  input      [7:0]    weights_payload_1_0_0_1,
  input      [7:0]    weights_payload_1_0_0_2,
  input      [7:0]    weights_payload_1_0_0_3,
  input      [7:0]    weights_payload_1_0_0_4,
  input      [7:0]    weights_payload_1_0_0_5,
  input      [7:0]    weights_payload_1_0_0_6,
  input      [7:0]    weights_payload_1_0_0_7,
  input      [7:0]    weights_payload_1_0_0_8,
  input      [7:0]    weights_payload_1_0_0_9,
  input      [7:0]    weights_payload_1_0_0_10,
  input      [7:0]    weights_payload_1_0_0_11,
  input      [7:0]    weights_payload_1_0_0_12,
  input      [7:0]    weights_payload_1_0_0_13,
  input      [7:0]    weights_payload_1_0_0_14,
  input      [7:0]    weights_payload_1_0_0_15,
  input      [7:0]    weights_payload_1_0_1_0,
  input      [7:0]    weights_payload_1_0_1_1,
  input      [7:0]    weights_payload_1_0_1_2,
  input      [7:0]    weights_payload_1_0_1_3,
  input      [7:0]    weights_payload_1_0_1_4,
  input      [7:0]    weights_payload_1_0_1_5,
  input      [7:0]    weights_payload_1_0_1_6,
  input      [7:0]    weights_payload_1_0_1_7,
  input      [7:0]    weights_payload_1_0_1_8,
  input      [7:0]    weights_payload_1_0_1_9,
  input      [7:0]    weights_payload_1_0_1_10,
  input      [7:0]    weights_payload_1_0_1_11,
  input      [7:0]    weights_payload_1_0_1_12,
  input      [7:0]    weights_payload_1_0_1_13,
  input      [7:0]    weights_payload_1_0_1_14,
  input      [7:0]    weights_payload_1_0_1_15,
  input      [7:0]    weights_payload_1_0_2_0,
  input      [7:0]    weights_payload_1_0_2_1,
  input      [7:0]    weights_payload_1_0_2_2,
  input      [7:0]    weights_payload_1_0_2_3,
  input      [7:0]    weights_payload_1_0_2_4,
  input      [7:0]    weights_payload_1_0_2_5,
  input      [7:0]    weights_payload_1_0_2_6,
  input      [7:0]    weights_payload_1_0_2_7,
  input      [7:0]    weights_payload_1_0_2_8,
  input      [7:0]    weights_payload_1_0_2_9,
  input      [7:0]    weights_payload_1_0_2_10,
  input      [7:0]    weights_payload_1_0_2_11,
  input      [7:0]    weights_payload_1_0_2_12,
  input      [7:0]    weights_payload_1_0_2_13,
  input      [7:0]    weights_payload_1_0_2_14,
  input      [7:0]    weights_payload_1_0_2_15,
  input      [7:0]    weights_payload_1_1_0_0,
  input      [7:0]    weights_payload_1_1_0_1,
  input      [7:0]    weights_payload_1_1_0_2,
  input      [7:0]    weights_payload_1_1_0_3,
  input      [7:0]    weights_payload_1_1_0_4,
  input      [7:0]    weights_payload_1_1_0_5,
  input      [7:0]    weights_payload_1_1_0_6,
  input      [7:0]    weights_payload_1_1_0_7,
  input      [7:0]    weights_payload_1_1_0_8,
  input      [7:0]    weights_payload_1_1_0_9,
  input      [7:0]    weights_payload_1_1_0_10,
  input      [7:0]    weights_payload_1_1_0_11,
  input      [7:0]    weights_payload_1_1_0_12,
  input      [7:0]    weights_payload_1_1_0_13,
  input      [7:0]    weights_payload_1_1_0_14,
  input      [7:0]    weights_payload_1_1_0_15,
  input      [7:0]    weights_payload_1_1_1_0,
  input      [7:0]    weights_payload_1_1_1_1,
  input      [7:0]    weights_payload_1_1_1_2,
  input      [7:0]    weights_payload_1_1_1_3,
  input      [7:0]    weights_payload_1_1_1_4,
  input      [7:0]    weights_payload_1_1_1_5,
  input      [7:0]    weights_payload_1_1_1_6,
  input      [7:0]    weights_payload_1_1_1_7,
  input      [7:0]    weights_payload_1_1_1_8,
  input      [7:0]    weights_payload_1_1_1_9,
  input      [7:0]    weights_payload_1_1_1_10,
  input      [7:0]    weights_payload_1_1_1_11,
  input      [7:0]    weights_payload_1_1_1_12,
  input      [7:0]    weights_payload_1_1_1_13,
  input      [7:0]    weights_payload_1_1_1_14,
  input      [7:0]    weights_payload_1_1_1_15,
  input      [7:0]    weights_payload_1_1_2_0,
  input      [7:0]    weights_payload_1_1_2_1,
  input      [7:0]    weights_payload_1_1_2_2,
  input      [7:0]    weights_payload_1_1_2_3,
  input      [7:0]    weights_payload_1_1_2_4,
  input      [7:0]    weights_payload_1_1_2_5,
  input      [7:0]    weights_payload_1_1_2_6,
  input      [7:0]    weights_payload_1_1_2_7,
  input      [7:0]    weights_payload_1_1_2_8,
  input      [7:0]    weights_payload_1_1_2_9,
  input      [7:0]    weights_payload_1_1_2_10,
  input      [7:0]    weights_payload_1_1_2_11,
  input      [7:0]    weights_payload_1_1_2_12,
  input      [7:0]    weights_payload_1_1_2_13,
  input      [7:0]    weights_payload_1_1_2_14,
  input      [7:0]    weights_payload_1_1_2_15,
  input      [7:0]    weights_payload_1_2_0_0,
  input      [7:0]    weights_payload_1_2_0_1,
  input      [7:0]    weights_payload_1_2_0_2,
  input      [7:0]    weights_payload_1_2_0_3,
  input      [7:0]    weights_payload_1_2_0_4,
  input      [7:0]    weights_payload_1_2_0_5,
  input      [7:0]    weights_payload_1_2_0_6,
  input      [7:0]    weights_payload_1_2_0_7,
  input      [7:0]    weights_payload_1_2_0_8,
  input      [7:0]    weights_payload_1_2_0_9,
  input      [7:0]    weights_payload_1_2_0_10,
  input      [7:0]    weights_payload_1_2_0_11,
  input      [7:0]    weights_payload_1_2_0_12,
  input      [7:0]    weights_payload_1_2_0_13,
  input      [7:0]    weights_payload_1_2_0_14,
  input      [7:0]    weights_payload_1_2_0_15,
  input      [7:0]    weights_payload_1_2_1_0,
  input      [7:0]    weights_payload_1_2_1_1,
  input      [7:0]    weights_payload_1_2_1_2,
  input      [7:0]    weights_payload_1_2_1_3,
  input      [7:0]    weights_payload_1_2_1_4,
  input      [7:0]    weights_payload_1_2_1_5,
  input      [7:0]    weights_payload_1_2_1_6,
  input      [7:0]    weights_payload_1_2_1_7,
  input      [7:0]    weights_payload_1_2_1_8,
  input      [7:0]    weights_payload_1_2_1_9,
  input      [7:0]    weights_payload_1_2_1_10,
  input      [7:0]    weights_payload_1_2_1_11,
  input      [7:0]    weights_payload_1_2_1_12,
  input      [7:0]    weights_payload_1_2_1_13,
  input      [7:0]    weights_payload_1_2_1_14,
  input      [7:0]    weights_payload_1_2_1_15,
  input      [7:0]    weights_payload_1_2_2_0,
  input      [7:0]    weights_payload_1_2_2_1,
  input      [7:0]    weights_payload_1_2_2_2,
  input      [7:0]    weights_payload_1_2_2_3,
  input      [7:0]    weights_payload_1_2_2_4,
  input      [7:0]    weights_payload_1_2_2_5,
  input      [7:0]    weights_payload_1_2_2_6,
  input      [7:0]    weights_payload_1_2_2_7,
  input      [7:0]    weights_payload_1_2_2_8,
  input      [7:0]    weights_payload_1_2_2_9,
  input      [7:0]    weights_payload_1_2_2_10,
  input      [7:0]    weights_payload_1_2_2_11,
  input      [7:0]    weights_payload_1_2_2_12,
  input      [7:0]    weights_payload_1_2_2_13,
  input      [7:0]    weights_payload_1_2_2_14,
  input      [7:0]    weights_payload_1_2_2_15,
  output              outputs_valid,
  input               outputs_ready,
  output     [23:0]   outputs_payload_frame_line_pixel_0,
  output     [23:0]   outputs_payload_frame_line_pixel_1,
  output              outputs_payload_frame_line_endOfLine,
  output              outputs_payload_frame_endOfFrame,
  output              outputs_payload_endOfPack,
  input               clk,
  input               reset
);

  wire                eventM2sPipes_9_eventIn_ready;
  wire                eventM2sPipes_9_eventOut_valid;
  wire                eventM2sPipes_9_CEs_0;
  wire                eventM2sPipes_9_CEs_1;
  wire                eventM2sPipes_9_CEs_2;
  wire                eventM2sPipes_9_CEs_3;
  wire                eventM2sPipes_9_CEs_4;
  wire                eventM2sPipes_9_CEs_5;
  wire                eventM2sPipes_9_CEs_6;
  wire                eventM2sPipes_9_CEs_7;
  wire                eventM2sPipes_9_CEs_8;
  wire       [15:0]   sIMD2INT8_1152_ab;
  wire       [15:0]   sIMD2INT8_1152_ac;
  wire       [15:0]   sIMD2INT8_1153_ab;
  wire       [15:0]   sIMD2INT8_1153_ac;
  wire       [15:0]   sIMD2INT8_1154_ab;
  wire       [15:0]   sIMD2INT8_1154_ac;
  wire       [15:0]   sIMD2INT8_1155_ab;
  wire       [15:0]   sIMD2INT8_1155_ac;
  wire       [15:0]   sIMD2INT8_1156_ab;
  wire       [15:0]   sIMD2INT8_1156_ac;
  wire       [15:0]   sIMD2INT8_1157_ab;
  wire       [15:0]   sIMD2INT8_1157_ac;
  wire       [15:0]   sIMD2INT8_1158_ab;
  wire       [15:0]   sIMD2INT8_1158_ac;
  wire       [15:0]   sIMD2INT8_1159_ab;
  wire       [15:0]   sIMD2INT8_1159_ac;
  wire       [15:0]   sIMD2INT8_1160_ab;
  wire       [15:0]   sIMD2INT8_1160_ac;
  wire       [15:0]   sIMD2INT8_1161_ab;
  wire       [15:0]   sIMD2INT8_1161_ac;
  wire       [15:0]   sIMD2INT8_1162_ab;
  wire       [15:0]   sIMD2INT8_1162_ac;
  wire       [15:0]   sIMD2INT8_1163_ab;
  wire       [15:0]   sIMD2INT8_1163_ac;
  wire       [15:0]   sIMD2INT8_1164_ab;
  wire       [15:0]   sIMD2INT8_1164_ac;
  wire       [15:0]   sIMD2INT8_1165_ab;
  wire       [15:0]   sIMD2INT8_1165_ac;
  wire       [15:0]   sIMD2INT8_1166_ab;
  wire       [15:0]   sIMD2INT8_1166_ac;
  wire       [15:0]   sIMD2INT8_1167_ab;
  wire       [15:0]   sIMD2INT8_1167_ac;
  wire       [15:0]   sIMD2INT8_1168_ab;
  wire       [15:0]   sIMD2INT8_1168_ac;
  wire       [15:0]   sIMD2INT8_1169_ab;
  wire       [15:0]   sIMD2INT8_1169_ac;
  wire       [15:0]   sIMD2INT8_1170_ab;
  wire       [15:0]   sIMD2INT8_1170_ac;
  wire       [15:0]   sIMD2INT8_1171_ab;
  wire       [15:0]   sIMD2INT8_1171_ac;
  wire       [15:0]   sIMD2INT8_1172_ab;
  wire       [15:0]   sIMD2INT8_1172_ac;
  wire       [15:0]   sIMD2INT8_1173_ab;
  wire       [15:0]   sIMD2INT8_1173_ac;
  wire       [15:0]   sIMD2INT8_1174_ab;
  wire       [15:0]   sIMD2INT8_1174_ac;
  wire       [15:0]   sIMD2INT8_1175_ab;
  wire       [15:0]   sIMD2INT8_1175_ac;
  wire       [15:0]   sIMD2INT8_1176_ab;
  wire       [15:0]   sIMD2INT8_1176_ac;
  wire       [15:0]   sIMD2INT8_1177_ab;
  wire       [15:0]   sIMD2INT8_1177_ac;
  wire       [15:0]   sIMD2INT8_1178_ab;
  wire       [15:0]   sIMD2INT8_1178_ac;
  wire       [15:0]   sIMD2INT8_1179_ab;
  wire       [15:0]   sIMD2INT8_1179_ac;
  wire       [15:0]   sIMD2INT8_1180_ab;
  wire       [15:0]   sIMD2INT8_1180_ac;
  wire       [15:0]   sIMD2INT8_1181_ab;
  wire       [15:0]   sIMD2INT8_1181_ac;
  wire       [15:0]   sIMD2INT8_1182_ab;
  wire       [15:0]   sIMD2INT8_1182_ac;
  wire       [15:0]   sIMD2INT8_1183_ab;
  wire       [15:0]   sIMD2INT8_1183_ac;
  wire       [15:0]   sIMD2INT8_1184_ab;
  wire       [15:0]   sIMD2INT8_1184_ac;
  wire       [15:0]   sIMD2INT8_1185_ab;
  wire       [15:0]   sIMD2INT8_1185_ac;
  wire       [15:0]   sIMD2INT8_1186_ab;
  wire       [15:0]   sIMD2INT8_1186_ac;
  wire       [15:0]   sIMD2INT8_1187_ab;
  wire       [15:0]   sIMD2INT8_1187_ac;
  wire       [15:0]   sIMD2INT8_1188_ab;
  wire       [15:0]   sIMD2INT8_1188_ac;
  wire       [15:0]   sIMD2INT8_1189_ab;
  wire       [15:0]   sIMD2INT8_1189_ac;
  wire       [15:0]   sIMD2INT8_1190_ab;
  wire       [15:0]   sIMD2INT8_1190_ac;
  wire       [15:0]   sIMD2INT8_1191_ab;
  wire       [15:0]   sIMD2INT8_1191_ac;
  wire       [15:0]   sIMD2INT8_1192_ab;
  wire       [15:0]   sIMD2INT8_1192_ac;
  wire       [15:0]   sIMD2INT8_1193_ab;
  wire       [15:0]   sIMD2INT8_1193_ac;
  wire       [15:0]   sIMD2INT8_1194_ab;
  wire       [15:0]   sIMD2INT8_1194_ac;
  wire       [15:0]   sIMD2INT8_1195_ab;
  wire       [15:0]   sIMD2INT8_1195_ac;
  wire       [15:0]   sIMD2INT8_1196_ab;
  wire       [15:0]   sIMD2INT8_1196_ac;
  wire       [15:0]   sIMD2INT8_1197_ab;
  wire       [15:0]   sIMD2INT8_1197_ac;
  wire       [15:0]   sIMD2INT8_1198_ab;
  wire       [15:0]   sIMD2INT8_1198_ac;
  wire       [15:0]   sIMD2INT8_1199_ab;
  wire       [15:0]   sIMD2INT8_1199_ac;
  wire       [15:0]   sIMD2INT8_1200_ab;
  wire       [15:0]   sIMD2INT8_1200_ac;
  wire       [15:0]   sIMD2INT8_1201_ab;
  wire       [15:0]   sIMD2INT8_1201_ac;
  wire       [15:0]   sIMD2INT8_1202_ab;
  wire       [15:0]   sIMD2INT8_1202_ac;
  wire       [15:0]   sIMD2INT8_1203_ab;
  wire       [15:0]   sIMD2INT8_1203_ac;
  wire       [15:0]   sIMD2INT8_1204_ab;
  wire       [15:0]   sIMD2INT8_1204_ac;
  wire       [15:0]   sIMD2INT8_1205_ab;
  wire       [15:0]   sIMD2INT8_1205_ac;
  wire       [15:0]   sIMD2INT8_1206_ab;
  wire       [15:0]   sIMD2INT8_1206_ac;
  wire       [15:0]   sIMD2INT8_1207_ab;
  wire       [15:0]   sIMD2INT8_1207_ac;
  wire       [15:0]   sIMD2INT8_1208_ab;
  wire       [15:0]   sIMD2INT8_1208_ac;
  wire       [15:0]   sIMD2INT8_1209_ab;
  wire       [15:0]   sIMD2INT8_1209_ac;
  wire       [15:0]   sIMD2INT8_1210_ab;
  wire       [15:0]   sIMD2INT8_1210_ac;
  wire       [15:0]   sIMD2INT8_1211_ab;
  wire       [15:0]   sIMD2INT8_1211_ac;
  wire       [15:0]   sIMD2INT8_1212_ab;
  wire       [15:0]   sIMD2INT8_1212_ac;
  wire       [15:0]   sIMD2INT8_1213_ab;
  wire       [15:0]   sIMD2INT8_1213_ac;
  wire       [15:0]   sIMD2INT8_1214_ab;
  wire       [15:0]   sIMD2INT8_1214_ac;
  wire       [15:0]   sIMD2INT8_1215_ab;
  wire       [15:0]   sIMD2INT8_1215_ac;
  wire       [15:0]   sIMD2INT8_1216_ab;
  wire       [15:0]   sIMD2INT8_1216_ac;
  wire       [15:0]   sIMD2INT8_1217_ab;
  wire       [15:0]   sIMD2INT8_1217_ac;
  wire       [15:0]   sIMD2INT8_1218_ab;
  wire       [15:0]   sIMD2INT8_1218_ac;
  wire       [15:0]   sIMD2INT8_1219_ab;
  wire       [15:0]   sIMD2INT8_1219_ac;
  wire       [15:0]   sIMD2INT8_1220_ab;
  wire       [15:0]   sIMD2INT8_1220_ac;
  wire       [15:0]   sIMD2INT8_1221_ab;
  wire       [15:0]   sIMD2INT8_1221_ac;
  wire       [15:0]   sIMD2INT8_1222_ab;
  wire       [15:0]   sIMD2INT8_1222_ac;
  wire       [15:0]   sIMD2INT8_1223_ab;
  wire       [15:0]   sIMD2INT8_1223_ac;
  wire       [15:0]   sIMD2INT8_1224_ab;
  wire       [15:0]   sIMD2INT8_1224_ac;
  wire       [15:0]   sIMD2INT8_1225_ab;
  wire       [15:0]   sIMD2INT8_1225_ac;
  wire       [15:0]   sIMD2INT8_1226_ab;
  wire       [15:0]   sIMD2INT8_1226_ac;
  wire       [15:0]   sIMD2INT8_1227_ab;
  wire       [15:0]   sIMD2INT8_1227_ac;
  wire       [15:0]   sIMD2INT8_1228_ab;
  wire       [15:0]   sIMD2INT8_1228_ac;
  wire       [15:0]   sIMD2INT8_1229_ab;
  wire       [15:0]   sIMD2INT8_1229_ac;
  wire       [15:0]   sIMD2INT8_1230_ab;
  wire       [15:0]   sIMD2INT8_1230_ac;
  wire       [15:0]   sIMD2INT8_1231_ab;
  wire       [15:0]   sIMD2INT8_1231_ac;
  wire       [15:0]   sIMD2INT8_1232_ab;
  wire       [15:0]   sIMD2INT8_1232_ac;
  wire       [15:0]   sIMD2INT8_1233_ab;
  wire       [15:0]   sIMD2INT8_1233_ac;
  wire       [15:0]   sIMD2INT8_1234_ab;
  wire       [15:0]   sIMD2INT8_1234_ac;
  wire       [15:0]   sIMD2INT8_1235_ab;
  wire       [15:0]   sIMD2INT8_1235_ac;
  wire       [15:0]   sIMD2INT8_1236_ab;
  wire       [15:0]   sIMD2INT8_1236_ac;
  wire       [15:0]   sIMD2INT8_1237_ab;
  wire       [15:0]   sIMD2INT8_1237_ac;
  wire       [15:0]   sIMD2INT8_1238_ab;
  wire       [15:0]   sIMD2INT8_1238_ac;
  wire       [15:0]   sIMD2INT8_1239_ab;
  wire       [15:0]   sIMD2INT8_1239_ac;
  wire       [15:0]   sIMD2INT8_1240_ab;
  wire       [15:0]   sIMD2INT8_1240_ac;
  wire       [15:0]   sIMD2INT8_1241_ab;
  wire       [15:0]   sIMD2INT8_1241_ac;
  wire       [15:0]   sIMD2INT8_1242_ab;
  wire       [15:0]   sIMD2INT8_1242_ac;
  wire       [15:0]   sIMD2INT8_1243_ab;
  wire       [15:0]   sIMD2INT8_1243_ac;
  wire       [15:0]   sIMD2INT8_1244_ab;
  wire       [15:0]   sIMD2INT8_1244_ac;
  wire       [15:0]   sIMD2INT8_1245_ab;
  wire       [15:0]   sIMD2INT8_1245_ac;
  wire       [15:0]   sIMD2INT8_1246_ab;
  wire       [15:0]   sIMD2INT8_1246_ac;
  wire       [15:0]   sIMD2INT8_1247_ab;
  wire       [15:0]   sIMD2INT8_1247_ac;
  wire       [15:0]   sIMD2INT8_1248_ab;
  wire       [15:0]   sIMD2INT8_1248_ac;
  wire       [15:0]   sIMD2INT8_1249_ab;
  wire       [15:0]   sIMD2INT8_1249_ac;
  wire       [15:0]   sIMD2INT8_1250_ab;
  wire       [15:0]   sIMD2INT8_1250_ac;
  wire       [15:0]   sIMD2INT8_1251_ab;
  wire       [15:0]   sIMD2INT8_1251_ac;
  wire       [15:0]   sIMD2INT8_1252_ab;
  wire       [15:0]   sIMD2INT8_1252_ac;
  wire       [15:0]   sIMD2INT8_1253_ab;
  wire       [15:0]   sIMD2INT8_1253_ac;
  wire       [15:0]   sIMD2INT8_1254_ab;
  wire       [15:0]   sIMD2INT8_1254_ac;
  wire       [15:0]   sIMD2INT8_1255_ab;
  wire       [15:0]   sIMD2INT8_1255_ac;
  wire       [15:0]   sIMD2INT8_1256_ab;
  wire       [15:0]   sIMD2INT8_1256_ac;
  wire       [15:0]   sIMD2INT8_1257_ab;
  wire       [15:0]   sIMD2INT8_1257_ac;
  wire       [15:0]   sIMD2INT8_1258_ab;
  wire       [15:0]   sIMD2INT8_1258_ac;
  wire       [15:0]   sIMD2INT8_1259_ab;
  wire       [15:0]   sIMD2INT8_1259_ac;
  wire       [15:0]   sIMD2INT8_1260_ab;
  wire       [15:0]   sIMD2INT8_1260_ac;
  wire       [15:0]   sIMD2INT8_1261_ab;
  wire       [15:0]   sIMD2INT8_1261_ac;
  wire       [15:0]   sIMD2INT8_1262_ab;
  wire       [15:0]   sIMD2INT8_1262_ac;
  wire       [15:0]   sIMD2INT8_1263_ab;
  wire       [15:0]   sIMD2INT8_1263_ac;
  wire       [15:0]   sIMD2INT8_1264_ab;
  wire       [15:0]   sIMD2INT8_1264_ac;
  wire       [15:0]   sIMD2INT8_1265_ab;
  wire       [15:0]   sIMD2INT8_1265_ac;
  wire       [15:0]   sIMD2INT8_1266_ab;
  wire       [15:0]   sIMD2INT8_1266_ac;
  wire       [15:0]   sIMD2INT8_1267_ab;
  wire       [15:0]   sIMD2INT8_1267_ac;
  wire       [15:0]   sIMD2INT8_1268_ab;
  wire       [15:0]   sIMD2INT8_1268_ac;
  wire       [15:0]   sIMD2INT8_1269_ab;
  wire       [15:0]   sIMD2INT8_1269_ac;
  wire       [15:0]   sIMD2INT8_1270_ab;
  wire       [15:0]   sIMD2INT8_1270_ac;
  wire       [15:0]   sIMD2INT8_1271_ab;
  wire       [15:0]   sIMD2INT8_1271_ac;
  wire       [15:0]   sIMD2INT8_1272_ab;
  wire       [15:0]   sIMD2INT8_1272_ac;
  wire       [15:0]   sIMD2INT8_1273_ab;
  wire       [15:0]   sIMD2INT8_1273_ac;
  wire       [15:0]   sIMD2INT8_1274_ab;
  wire       [15:0]   sIMD2INT8_1274_ac;
  wire       [15:0]   sIMD2INT8_1275_ab;
  wire       [15:0]   sIMD2INT8_1275_ac;
  wire       [15:0]   sIMD2INT8_1276_ab;
  wire       [15:0]   sIMD2INT8_1276_ac;
  wire       [15:0]   sIMD2INT8_1277_ab;
  wire       [15:0]   sIMD2INT8_1277_ac;
  wire       [15:0]   sIMD2INT8_1278_ab;
  wire       [15:0]   sIMD2INT8_1278_ac;
  wire       [15:0]   sIMD2INT8_1279_ab;
  wire       [15:0]   sIMD2INT8_1279_ac;
  wire       [15:0]   sIMD2INT8_1280_ab;
  wire       [15:0]   sIMD2INT8_1280_ac;
  wire       [15:0]   sIMD2INT8_1281_ab;
  wire       [15:0]   sIMD2INT8_1281_ac;
  wire       [15:0]   sIMD2INT8_1282_ab;
  wire       [15:0]   sIMD2INT8_1282_ac;
  wire       [15:0]   sIMD2INT8_1283_ab;
  wire       [15:0]   sIMD2INT8_1283_ac;
  wire       [15:0]   sIMD2INT8_1284_ab;
  wire       [15:0]   sIMD2INT8_1284_ac;
  wire       [15:0]   sIMD2INT8_1285_ab;
  wire       [15:0]   sIMD2INT8_1285_ac;
  wire       [15:0]   sIMD2INT8_1286_ab;
  wire       [15:0]   sIMD2INT8_1286_ac;
  wire       [15:0]   sIMD2INT8_1287_ab;
  wire       [15:0]   sIMD2INT8_1287_ac;
  wire       [15:0]   sIMD2INT8_1288_ab;
  wire       [15:0]   sIMD2INT8_1288_ac;
  wire       [15:0]   sIMD2INT8_1289_ab;
  wire       [15:0]   sIMD2INT8_1289_ac;
  wire       [15:0]   sIMD2INT8_1290_ab;
  wire       [15:0]   sIMD2INT8_1290_ac;
  wire       [15:0]   sIMD2INT8_1291_ab;
  wire       [15:0]   sIMD2INT8_1291_ac;
  wire       [15:0]   sIMD2INT8_1292_ab;
  wire       [15:0]   sIMD2INT8_1292_ac;
  wire       [15:0]   sIMD2INT8_1293_ab;
  wire       [15:0]   sIMD2INT8_1293_ac;
  wire       [15:0]   sIMD2INT8_1294_ab;
  wire       [15:0]   sIMD2INT8_1294_ac;
  wire       [15:0]   sIMD2INT8_1295_ab;
  wire       [15:0]   sIMD2INT8_1295_ac;
  wire                acc_videoIn_ready;
  wire                acc_videoOut_valid;
  wire       [23:0]   acc_videoOut_payload_frame_line_pixel_0;
  wire       [23:0]   acc_videoOut_payload_frame_line_pixel_1;
  wire                acc_videoOut_payload_frame_line_endOfLine;
  wire                acc_videoOut_payload_frame_endOfFrame;
  wire                acc_videoOut_payload_endOfPack;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_1;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_2;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_3;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_4;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_5;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_6;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_7;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_8;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_9;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_10;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_11;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_12;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_13;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_14;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_15;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_16;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_17;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_18;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_19;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_20;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_21;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_22;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_23;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_24;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_25;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_26;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_27;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_28;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_29;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_30;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_31;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_32;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_33;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_34;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_35;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_36;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_37;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_38;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_39;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_40;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_41;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_42;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_43;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_44;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_45;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_46;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_47;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_48;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_49;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_50;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_51;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_52;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_53;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_54;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_55;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_56;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_57;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_58;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_59;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_60;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_61;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_62;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_63;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_64;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_65;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_66;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_67;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_68;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_70;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_71;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_72;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_0_72_1;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_1;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_2;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_3;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_4;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_5;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_6;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_7;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_8;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_9;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_10;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_11;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_12;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_13;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_14;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_15;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_16;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_17;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_18;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_19;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_20;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_21;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_22;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_23;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_24;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_25;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_26;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_27;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_28;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_29;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_30;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_31;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_32;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_33;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_34;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_35;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_36;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_37;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_38;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_39;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_40;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_41;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_42;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_43;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_44;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_45;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_46;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_47;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_48;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_49;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_50;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_51;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_52;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_53;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_54;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_55;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_56;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_57;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_58;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_59;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_60;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_61;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_62;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_63;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_64;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_65;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_66;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_67;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_68;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_70;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_71;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_72;
  wire       [15:0]   tmp_tmp_postConv_payload_frame_line_pixel_1_72_1;
  wire                tmp_inputs_ready;
  wire                inputsT_valid;
  wire                inputsT_ready;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    inputsT_payload_frame_line_pixel_2_2_15;
  wire                inputsT_payload_frame_line_endOfLine;
  wire                inputsT_payload_frame_endOfFrame;
  wire                inputsT_payload_endOfPack;
  wire                prevConv_valid;
  wire                prevConv_ready;
  wire       [7:0]    prevConv_payload_frame_line_pixel_0_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_0_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_0_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_1_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_1_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_1_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_2_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_2_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_2_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_3_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_3_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_3_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_4_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_4_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_4_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_5_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_5_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_5_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_6_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_6_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_6_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_7_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_7_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_7_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_8_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_8_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_8_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_9_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_9_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_9_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_10_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_10_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_10_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_11_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_11_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_11_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_12_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_12_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_12_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_13_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_13_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_13_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_14_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_14_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_14_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_15_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_15_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_15_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_16_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_16_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_16_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_17_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_17_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_17_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_18_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_18_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_18_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_19_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_19_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_19_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_20_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_20_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_20_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_21_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_21_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_21_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_22_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_22_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_22_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_23_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_23_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_23_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_24_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_24_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_24_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_25_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_25_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_25_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_26_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_26_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_26_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_27_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_27_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_27_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_28_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_28_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_28_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_29_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_29_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_29_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_30_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_30_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_30_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_31_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_31_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_31_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_32_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_32_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_32_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_33_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_33_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_33_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_34_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_34_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_34_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_35_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_35_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_35_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_36_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_36_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_36_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_37_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_37_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_37_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_38_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_38_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_38_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_39_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_39_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_39_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_40_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_40_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_40_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_41_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_41_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_41_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_42_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_42_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_42_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_43_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_43_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_43_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_44_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_44_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_44_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_45_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_45_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_45_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_46_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_46_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_46_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_47_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_47_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_47_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_48_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_48_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_48_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_49_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_49_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_49_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_50_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_50_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_50_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_51_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_51_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_51_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_52_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_52_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_52_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_53_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_53_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_53_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_54_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_54_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_54_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_55_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_55_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_55_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_56_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_56_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_56_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_57_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_57_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_57_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_58_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_58_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_58_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_59_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_59_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_59_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_60_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_60_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_60_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_61_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_61_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_61_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_62_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_62_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_62_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_63_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_63_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_63_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_64_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_64_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_64_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_65_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_65_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_65_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_66_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_66_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_66_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_67_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_67_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_67_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_68_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_68_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_68_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_69_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_69_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_69_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_70_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_70_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_70_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_71_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_71_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_71_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_72_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_72_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_72_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_73_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_73_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_73_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_74_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_74_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_74_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_75_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_75_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_75_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_76_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_76_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_76_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_77_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_77_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_77_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_78_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_78_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_78_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_79_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_79_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_79_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_80_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_80_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_80_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_81_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_81_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_81_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_82_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_82_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_82_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_83_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_83_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_83_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_84_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_84_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_84_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_85_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_85_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_85_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_86_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_86_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_86_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_87_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_87_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_87_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_88_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_88_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_88_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_89_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_89_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_89_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_90_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_90_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_90_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_91_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_91_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_91_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_92_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_92_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_92_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_93_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_93_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_93_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_94_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_94_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_94_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_95_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_95_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_95_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_96_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_96_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_96_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_97_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_97_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_97_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_98_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_98_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_98_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_99_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_99_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_99_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_100_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_100_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_100_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_101_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_101_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_101_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_102_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_102_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_102_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_103_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_103_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_103_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_104_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_104_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_104_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_105_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_105_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_105_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_106_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_106_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_106_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_107_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_107_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_107_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_108_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_108_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_108_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_109_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_109_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_109_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_110_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_110_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_110_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_111_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_111_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_111_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_112_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_112_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_112_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_113_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_113_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_113_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_114_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_114_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_114_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_115_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_115_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_115_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_116_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_116_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_116_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_117_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_117_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_117_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_118_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_118_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_118_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_119_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_119_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_119_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_120_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_120_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_120_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_121_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_121_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_121_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_122_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_122_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_122_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_123_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_123_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_123_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_124_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_124_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_124_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_125_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_125_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_125_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_126_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_126_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_126_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_127_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_127_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_127_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_128_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_128_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_128_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_129_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_129_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_129_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_130_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_130_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_130_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_131_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_131_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_131_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_132_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_132_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_132_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_133_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_133_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_133_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_134_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_134_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_134_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_135_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_135_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_135_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_136_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_136_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_136_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_137_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_137_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_137_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_138_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_138_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_138_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_139_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_139_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_139_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_140_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_140_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_140_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_141_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_141_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_141_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_142_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_142_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_142_2;
  wire       [7:0]    prevConv_payload_frame_line_pixel_143_0;
  wire       [7:0]    prevConv_payload_frame_line_pixel_143_1;
  wire       [7:0]    prevConv_payload_frame_line_pixel_143_2;
  wire                prevConv_payload_frame_line_endOfLine;
  wire                prevConv_payload_frame_endOfFrame;
  wire                prevConv_payload_endOfPack;
  wire                postConv_valid;
  wire                postConv_ready;
  wire       [15:0]   postConv_payload_frame_line_pixel_0;
  wire       [15:0]   postConv_payload_frame_line_pixel_1;
  wire                postConv_payload_frame_line_endOfLine;
  wire                postConv_payload_frame_endOfFrame;
  wire                postConv_payload_endOfPack;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_1;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_2;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_3;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_4;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_5;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_6;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_7;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_8;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_9;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_10;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_11;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_12;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_13;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_14;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_15;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_16;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_17;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_18;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_19;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_20;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_21;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_22;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_23;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_24;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_25;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_26;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_27;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_28;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_29;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_30;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_31;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_32;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_33;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_34;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_35;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_36;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_37;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_38;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_39;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_40;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_41;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_42;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_43;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_44;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_45;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_46;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_47;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_48;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_49;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_50;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_51;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_52;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_53;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_54;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_55;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_56;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_57;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_58;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_59;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_60;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_61;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_62;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_63;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_64;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_65;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_66;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_67;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_68;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_69;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_70;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_71;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_0_72;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_1;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_2;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_3;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_4;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_5;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_6;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_7;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_8;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_9;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_10;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_11;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_12;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_13;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_14;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_15;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_16;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_17;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_18;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_19;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_20;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_21;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_22;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_23;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_24;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_25;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_26;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_27;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_28;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_29;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_30;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_31;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_32;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_33;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_34;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_35;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_36;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_37;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_38;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_39;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_40;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_41;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_42;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_43;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_44;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_45;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_46;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_47;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_48;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_49;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_50;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_51;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_52;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_53;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_54;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_55;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_56;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_57;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_58;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_59;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_60;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_61;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_62;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_63;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_64;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_65;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_66;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_67;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_68;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_69;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_70;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_71;
  reg        [15:0]   tmp_postConv_payload_frame_line_pixel_1_72;
  reg                 tmp_postConv_payload_frame_line_endOfLine;
  reg                 tmp_postConv_payload_frame_endOfFrame;
  reg                 tmp_postConv_payload_endOfPack;
  reg                 tmp_postConv_payload_frame_line_endOfLine_1;
  reg                 tmp_postConv_payload_frame_endOfFrame_1;
  reg                 tmp_postConv_payload_endOfPack_1;
  reg                 tmp_postConv_payload_frame_line_endOfLine_2;
  reg                 tmp_postConv_payload_frame_endOfFrame_2;
  reg                 tmp_postConv_payload_endOfPack_2;
  reg                 tmp_postConv_payload_frame_line_endOfLine_3;
  reg                 tmp_postConv_payload_frame_endOfFrame_3;
  reg                 tmp_postConv_payload_endOfPack_3;
  reg                 tmp_postConv_payload_frame_line_endOfLine_4;
  reg                 tmp_postConv_payload_frame_endOfFrame_4;
  reg                 tmp_postConv_payload_endOfPack_4;
  reg                 tmp_postConv_payload_frame_line_endOfLine_5;
  reg                 tmp_postConv_payload_frame_endOfFrame_5;
  reg                 tmp_postConv_payload_endOfPack_5;
  reg                 tmp_postConv_payload_frame_line_endOfLine_6;
  reg                 tmp_postConv_payload_frame_endOfFrame_6;
  reg                 tmp_postConv_payload_endOfPack_6;
  reg                 tmp_postConv_payload_frame_line_endOfLine_7;
  reg                 tmp_postConv_payload_frame_endOfFrame_7;
  reg                 tmp_postConv_payload_endOfPack_7;
  reg                 tmp_postConv_payload_frame_line_endOfLine_8;
  reg                 tmp_postConv_payload_frame_endOfFrame_8;
  reg                 tmp_postConv_payload_endOfPack_8;
  wire                inputsT_fire;
  wire                postConv_s2mPipe_valid;
  wire                postConv_s2mPipe_ready;
  wire       [15:0]   postConv_s2mPipe_payload_frame_line_pixel_0;
  wire       [15:0]   postConv_s2mPipe_payload_frame_line_pixel_1;
  wire                postConv_s2mPipe_payload_frame_line_endOfLine;
  wire                postConv_s2mPipe_payload_frame_endOfFrame;
  wire                postConv_s2mPipe_payload_endOfPack;
  reg                 postConv_rValid;
  reg        [15:0]   postConv_rData_frame_line_pixel_0;
  reg        [15:0]   postConv_rData_frame_line_pixel_1;
  reg                 postConv_rData_frame_line_endOfLine;
  reg                 postConv_rData_frame_endOfFrame;
  reg                 postConv_rData_endOfPack;

  assign tmp_tmp_postConv_payload_frame_line_pixel_0 = ($signed(sIMD2INT8_1152_ab) + $signed(sIMD2INT8_1153_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_1 = ($signed(sIMD2INT8_1155_ab) + $signed(sIMD2INT8_1156_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_2 = ($signed(sIMD2INT8_1158_ab) + $signed(sIMD2INT8_1159_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_3 = ($signed(sIMD2INT8_1161_ab) + $signed(sIMD2INT8_1162_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_4 = ($signed(sIMD2INT8_1164_ab) + $signed(sIMD2INT8_1165_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_5 = ($signed(sIMD2INT8_1167_ab) + $signed(sIMD2INT8_1168_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_6 = ($signed(sIMD2INT8_1170_ab) + $signed(sIMD2INT8_1171_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_7 = ($signed(sIMD2INT8_1173_ab) + $signed(sIMD2INT8_1174_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_8 = ($signed(sIMD2INT8_1176_ab) + $signed(sIMD2INT8_1177_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_9 = ($signed(sIMD2INT8_1179_ab) + $signed(sIMD2INT8_1180_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_10 = ($signed(sIMD2INT8_1182_ab) + $signed(sIMD2INT8_1183_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_11 = ($signed(sIMD2INT8_1185_ab) + $signed(sIMD2INT8_1186_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_12 = ($signed(sIMD2INT8_1188_ab) + $signed(sIMD2INT8_1189_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_13 = ($signed(sIMD2INT8_1191_ab) + $signed(sIMD2INT8_1192_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_14 = ($signed(sIMD2INT8_1194_ab) + $signed(sIMD2INT8_1195_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_15 = ($signed(sIMD2INT8_1197_ab) + $signed(sIMD2INT8_1198_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_16 = ($signed(sIMD2INT8_1200_ab) + $signed(sIMD2INT8_1201_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_17 = ($signed(sIMD2INT8_1203_ab) + $signed(sIMD2INT8_1204_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_18 = ($signed(sIMD2INT8_1206_ab) + $signed(sIMD2INT8_1207_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_19 = ($signed(sIMD2INT8_1209_ab) + $signed(sIMD2INT8_1210_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_20 = ($signed(sIMD2INT8_1212_ab) + $signed(sIMD2INT8_1213_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_21 = ($signed(sIMD2INT8_1215_ab) + $signed(sIMD2INT8_1216_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_22 = ($signed(sIMD2INT8_1218_ab) + $signed(sIMD2INT8_1219_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_23 = ($signed(sIMD2INT8_1221_ab) + $signed(sIMD2INT8_1222_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_24 = ($signed(sIMD2INT8_1224_ab) + $signed(sIMD2INT8_1225_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_25 = ($signed(sIMD2INT8_1227_ab) + $signed(sIMD2INT8_1228_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_26 = ($signed(sIMD2INT8_1230_ab) + $signed(sIMD2INT8_1231_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_27 = ($signed(sIMD2INT8_1233_ab) + $signed(sIMD2INT8_1234_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_28 = ($signed(sIMD2INT8_1236_ab) + $signed(sIMD2INT8_1237_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_29 = ($signed(sIMD2INT8_1239_ab) + $signed(sIMD2INT8_1240_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_30 = ($signed(sIMD2INT8_1242_ab) + $signed(sIMD2INT8_1243_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_31 = ($signed(sIMD2INT8_1245_ab) + $signed(sIMD2INT8_1246_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_32 = ($signed(sIMD2INT8_1248_ab) + $signed(sIMD2INT8_1249_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_33 = ($signed(sIMD2INT8_1251_ab) + $signed(sIMD2INT8_1252_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_34 = ($signed(sIMD2INT8_1254_ab) + $signed(sIMD2INT8_1255_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_35 = ($signed(sIMD2INT8_1257_ab) + $signed(sIMD2INT8_1258_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_36 = ($signed(sIMD2INT8_1260_ab) + $signed(sIMD2INT8_1261_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_37 = ($signed(sIMD2INT8_1263_ab) + $signed(sIMD2INT8_1264_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_38 = ($signed(sIMD2INT8_1266_ab) + $signed(sIMD2INT8_1267_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_39 = ($signed(sIMD2INT8_1269_ab) + $signed(sIMD2INT8_1270_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_40 = ($signed(sIMD2INT8_1272_ab) + $signed(sIMD2INT8_1273_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_41 = ($signed(sIMD2INT8_1275_ab) + $signed(sIMD2INT8_1276_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_42 = ($signed(sIMD2INT8_1278_ab) + $signed(sIMD2INT8_1279_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_43 = ($signed(sIMD2INT8_1281_ab) + $signed(sIMD2INT8_1282_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_44 = ($signed(sIMD2INT8_1284_ab) + $signed(sIMD2INT8_1285_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_45 = ($signed(sIMD2INT8_1287_ab) + $signed(sIMD2INT8_1288_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_46 = ($signed(sIMD2INT8_1290_ab) + $signed(sIMD2INT8_1291_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_47 = ($signed(sIMD2INT8_1293_ab) + $signed(sIMD2INT8_1294_ab));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_48 = ($signed(tmp_postConv_payload_frame_line_pixel_0) + $signed(tmp_postConv_payload_frame_line_pixel_0_1));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_49 = ($signed(tmp_postConv_payload_frame_line_pixel_0_3) + $signed(tmp_postConv_payload_frame_line_pixel_0_4));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_50 = ($signed(tmp_postConv_payload_frame_line_pixel_0_6) + $signed(tmp_postConv_payload_frame_line_pixel_0_7));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_51 = ($signed(tmp_postConv_payload_frame_line_pixel_0_9) + $signed(tmp_postConv_payload_frame_line_pixel_0_10));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_52 = ($signed(tmp_postConv_payload_frame_line_pixel_0_12) + $signed(tmp_postConv_payload_frame_line_pixel_0_13));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_53 = ($signed(tmp_postConv_payload_frame_line_pixel_0_15) + $signed(tmp_postConv_payload_frame_line_pixel_0_16));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_54 = ($signed(tmp_postConv_payload_frame_line_pixel_0_18) + $signed(tmp_postConv_payload_frame_line_pixel_0_19));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_55 = ($signed(tmp_postConv_payload_frame_line_pixel_0_21) + $signed(tmp_postConv_payload_frame_line_pixel_0_22));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_56 = ($signed(tmp_postConv_payload_frame_line_pixel_0_24) + $signed(tmp_postConv_payload_frame_line_pixel_0_25));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_57 = ($signed(tmp_postConv_payload_frame_line_pixel_0_27) + $signed(tmp_postConv_payload_frame_line_pixel_0_28));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_58 = ($signed(tmp_postConv_payload_frame_line_pixel_0_30) + $signed(tmp_postConv_payload_frame_line_pixel_0_31));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_59 = ($signed(tmp_postConv_payload_frame_line_pixel_0_33) + $signed(tmp_postConv_payload_frame_line_pixel_0_34));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_60 = ($signed(tmp_postConv_payload_frame_line_pixel_0_36) + $signed(tmp_postConv_payload_frame_line_pixel_0_37));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_61 = ($signed(tmp_postConv_payload_frame_line_pixel_0_39) + $signed(tmp_postConv_payload_frame_line_pixel_0_40));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_62 = ($signed(tmp_postConv_payload_frame_line_pixel_0_42) + $signed(tmp_postConv_payload_frame_line_pixel_0_43));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_63 = ($signed(tmp_postConv_payload_frame_line_pixel_0_45) + $signed(tmp_postConv_payload_frame_line_pixel_0_46));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_64 = ($signed(tmp_postConv_payload_frame_line_pixel_0_48) + $signed(tmp_postConv_payload_frame_line_pixel_0_49));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_65 = ($signed(tmp_postConv_payload_frame_line_pixel_0_51) + $signed(tmp_postConv_payload_frame_line_pixel_0_52));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_66 = ($signed(tmp_postConv_payload_frame_line_pixel_0_54) + $signed(tmp_postConv_payload_frame_line_pixel_0_55));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_67 = ($signed(tmp_postConv_payload_frame_line_pixel_0_57) + $signed(tmp_postConv_payload_frame_line_pixel_0_58));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_68 = ($signed(tmp_postConv_payload_frame_line_pixel_0_60) + $signed(tmp_postConv_payload_frame_line_pixel_0_61));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_70 = ($signed(tmp_postConv_payload_frame_line_pixel_0_64) + $signed(tmp_postConv_payload_frame_line_pixel_0_65));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_71 = ($signed(tmp_postConv_payload_frame_line_pixel_0_67) + $signed(tmp_postConv_payload_frame_line_pixel_0_68));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_72 = ($signed(tmp_postConv_payload_frame_line_pixel_0_70) + $signed(tmp_postConv_payload_frame_line_pixel_0_71));
  assign tmp_tmp_postConv_payload_frame_line_pixel_0_72_1 = 16'h0;
  assign tmp_tmp_postConv_payload_frame_line_pixel_1 = ($signed(sIMD2INT8_1152_ac) + $signed(sIMD2INT8_1153_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_1 = ($signed(sIMD2INT8_1155_ac) + $signed(sIMD2INT8_1156_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_2 = ($signed(sIMD2INT8_1158_ac) + $signed(sIMD2INT8_1159_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_3 = ($signed(sIMD2INT8_1161_ac) + $signed(sIMD2INT8_1162_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_4 = ($signed(sIMD2INT8_1164_ac) + $signed(sIMD2INT8_1165_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_5 = ($signed(sIMD2INT8_1167_ac) + $signed(sIMD2INT8_1168_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_6 = ($signed(sIMD2INT8_1170_ac) + $signed(sIMD2INT8_1171_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_7 = ($signed(sIMD2INT8_1173_ac) + $signed(sIMD2INT8_1174_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_8 = ($signed(sIMD2INT8_1176_ac) + $signed(sIMD2INT8_1177_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_9 = ($signed(sIMD2INT8_1179_ac) + $signed(sIMD2INT8_1180_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_10 = ($signed(sIMD2INT8_1182_ac) + $signed(sIMD2INT8_1183_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_11 = ($signed(sIMD2INT8_1185_ac) + $signed(sIMD2INT8_1186_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_12 = ($signed(sIMD2INT8_1188_ac) + $signed(sIMD2INT8_1189_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_13 = ($signed(sIMD2INT8_1191_ac) + $signed(sIMD2INT8_1192_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_14 = ($signed(sIMD2INT8_1194_ac) + $signed(sIMD2INT8_1195_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_15 = ($signed(sIMD2INT8_1197_ac) + $signed(sIMD2INT8_1198_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_16 = ($signed(sIMD2INT8_1200_ac) + $signed(sIMD2INT8_1201_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_17 = ($signed(sIMD2INT8_1203_ac) + $signed(sIMD2INT8_1204_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_18 = ($signed(sIMD2INT8_1206_ac) + $signed(sIMD2INT8_1207_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_19 = ($signed(sIMD2INT8_1209_ac) + $signed(sIMD2INT8_1210_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_20 = ($signed(sIMD2INT8_1212_ac) + $signed(sIMD2INT8_1213_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_21 = ($signed(sIMD2INT8_1215_ac) + $signed(sIMD2INT8_1216_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_22 = ($signed(sIMD2INT8_1218_ac) + $signed(sIMD2INT8_1219_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_23 = ($signed(sIMD2INT8_1221_ac) + $signed(sIMD2INT8_1222_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_24 = ($signed(sIMD2INT8_1224_ac) + $signed(sIMD2INT8_1225_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_25 = ($signed(sIMD2INT8_1227_ac) + $signed(sIMD2INT8_1228_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_26 = ($signed(sIMD2INT8_1230_ac) + $signed(sIMD2INT8_1231_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_27 = ($signed(sIMD2INT8_1233_ac) + $signed(sIMD2INT8_1234_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_28 = ($signed(sIMD2INT8_1236_ac) + $signed(sIMD2INT8_1237_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_29 = ($signed(sIMD2INT8_1239_ac) + $signed(sIMD2INT8_1240_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_30 = ($signed(sIMD2INT8_1242_ac) + $signed(sIMD2INT8_1243_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_31 = ($signed(sIMD2INT8_1245_ac) + $signed(sIMD2INT8_1246_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_32 = ($signed(sIMD2INT8_1248_ac) + $signed(sIMD2INT8_1249_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_33 = ($signed(sIMD2INT8_1251_ac) + $signed(sIMD2INT8_1252_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_34 = ($signed(sIMD2INT8_1254_ac) + $signed(sIMD2INT8_1255_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_35 = ($signed(sIMD2INT8_1257_ac) + $signed(sIMD2INT8_1258_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_36 = ($signed(sIMD2INT8_1260_ac) + $signed(sIMD2INT8_1261_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_37 = ($signed(sIMD2INT8_1263_ac) + $signed(sIMD2INT8_1264_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_38 = ($signed(sIMD2INT8_1266_ac) + $signed(sIMD2INT8_1267_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_39 = ($signed(sIMD2INT8_1269_ac) + $signed(sIMD2INT8_1270_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_40 = ($signed(sIMD2INT8_1272_ac) + $signed(sIMD2INT8_1273_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_41 = ($signed(sIMD2INT8_1275_ac) + $signed(sIMD2INT8_1276_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_42 = ($signed(sIMD2INT8_1278_ac) + $signed(sIMD2INT8_1279_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_43 = ($signed(sIMD2INT8_1281_ac) + $signed(sIMD2INT8_1282_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_44 = ($signed(sIMD2INT8_1284_ac) + $signed(sIMD2INT8_1285_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_45 = ($signed(sIMD2INT8_1287_ac) + $signed(sIMD2INT8_1288_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_46 = ($signed(sIMD2INT8_1290_ac) + $signed(sIMD2INT8_1291_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_47 = ($signed(sIMD2INT8_1293_ac) + $signed(sIMD2INT8_1294_ac));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_48 = ($signed(tmp_postConv_payload_frame_line_pixel_1) + $signed(tmp_postConv_payload_frame_line_pixel_1_1));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_49 = ($signed(tmp_postConv_payload_frame_line_pixel_1_3) + $signed(tmp_postConv_payload_frame_line_pixel_1_4));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_50 = ($signed(tmp_postConv_payload_frame_line_pixel_1_6) + $signed(tmp_postConv_payload_frame_line_pixel_1_7));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_51 = ($signed(tmp_postConv_payload_frame_line_pixel_1_9) + $signed(tmp_postConv_payload_frame_line_pixel_1_10));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_52 = ($signed(tmp_postConv_payload_frame_line_pixel_1_12) + $signed(tmp_postConv_payload_frame_line_pixel_1_13));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_53 = ($signed(tmp_postConv_payload_frame_line_pixel_1_15) + $signed(tmp_postConv_payload_frame_line_pixel_1_16));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_54 = ($signed(tmp_postConv_payload_frame_line_pixel_1_18) + $signed(tmp_postConv_payload_frame_line_pixel_1_19));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_55 = ($signed(tmp_postConv_payload_frame_line_pixel_1_21) + $signed(tmp_postConv_payload_frame_line_pixel_1_22));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_56 = ($signed(tmp_postConv_payload_frame_line_pixel_1_24) + $signed(tmp_postConv_payload_frame_line_pixel_1_25));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_57 = ($signed(tmp_postConv_payload_frame_line_pixel_1_27) + $signed(tmp_postConv_payload_frame_line_pixel_1_28));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_58 = ($signed(tmp_postConv_payload_frame_line_pixel_1_30) + $signed(tmp_postConv_payload_frame_line_pixel_1_31));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_59 = ($signed(tmp_postConv_payload_frame_line_pixel_1_33) + $signed(tmp_postConv_payload_frame_line_pixel_1_34));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_60 = ($signed(tmp_postConv_payload_frame_line_pixel_1_36) + $signed(tmp_postConv_payload_frame_line_pixel_1_37));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_61 = ($signed(tmp_postConv_payload_frame_line_pixel_1_39) + $signed(tmp_postConv_payload_frame_line_pixel_1_40));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_62 = ($signed(tmp_postConv_payload_frame_line_pixel_1_42) + $signed(tmp_postConv_payload_frame_line_pixel_1_43));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_63 = ($signed(tmp_postConv_payload_frame_line_pixel_1_45) + $signed(tmp_postConv_payload_frame_line_pixel_1_46));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_64 = ($signed(tmp_postConv_payload_frame_line_pixel_1_48) + $signed(tmp_postConv_payload_frame_line_pixel_1_49));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_65 = ($signed(tmp_postConv_payload_frame_line_pixel_1_51) + $signed(tmp_postConv_payload_frame_line_pixel_1_52));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_66 = ($signed(tmp_postConv_payload_frame_line_pixel_1_54) + $signed(tmp_postConv_payload_frame_line_pixel_1_55));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_67 = ($signed(tmp_postConv_payload_frame_line_pixel_1_57) + $signed(tmp_postConv_payload_frame_line_pixel_1_58));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_68 = ($signed(tmp_postConv_payload_frame_line_pixel_1_60) + $signed(tmp_postConv_payload_frame_line_pixel_1_61));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_70 = ($signed(tmp_postConv_payload_frame_line_pixel_1_64) + $signed(tmp_postConv_payload_frame_line_pixel_1_65));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_71 = ($signed(tmp_postConv_payload_frame_line_pixel_1_67) + $signed(tmp_postConv_payload_frame_line_pixel_1_68));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_72 = ($signed(tmp_postConv_payload_frame_line_pixel_1_70) + $signed(tmp_postConv_payload_frame_line_pixel_1_71));
  assign tmp_tmp_postConv_payload_frame_line_pixel_1_72_1 = 16'h0;
  EventM2sPipes eventM2sPipes_9 (
    .eventIn_valid     (prevConv_valid                  ), //i
    .eventIn_ready     (eventM2sPipes_9_eventIn_ready   ), //o
    .eventOut_valid    (eventM2sPipes_9_eventOut_valid  ), //o
    .eventOut_ready    (postConv_ready                  ), //i
    .CEs_0             (eventM2sPipes_9_CEs_0           ), //o
    .CEs_1             (eventM2sPipes_9_CEs_1           ), //o
    .CEs_2             (eventM2sPipes_9_CEs_2           ), //o
    .CEs_3             (eventM2sPipes_9_CEs_3           ), //o
    .CEs_4             (eventM2sPipes_9_CEs_4           ), //o
    .CEs_5             (eventM2sPipes_9_CEs_5           ), //o
    .CEs_6             (eventM2sPipes_9_CEs_6           ), //o
    .CEs_7             (eventM2sPipes_9_CEs_7           ), //o
    .CEs_8             (eventM2sPipes_9_CEs_8           ), //o
    .clk               (clk                             ), //i
    .reset             (reset                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1152 (
    .a        (prevConv_payload_frame_line_pixel_0_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_0_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_0_2[7:0]  ), //i
    .ab       (sIMD2INT8_1152_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1152_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1153 (
    .a        (prevConv_payload_frame_line_pixel_1_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_1_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_1_2[7:0]  ), //i
    .ab       (sIMD2INT8_1153_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1153_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1154 (
    .a        (prevConv_payload_frame_line_pixel_2_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_2_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_2_2[7:0]  ), //i
    .ab       (sIMD2INT8_1154_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1154_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1155 (
    .a        (prevConv_payload_frame_line_pixel_3_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_3_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_3_2[7:0]  ), //i
    .ab       (sIMD2INT8_1155_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1155_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1156 (
    .a        (prevConv_payload_frame_line_pixel_4_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_4_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_4_2[7:0]  ), //i
    .ab       (sIMD2INT8_1156_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1156_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1157 (
    .a        (prevConv_payload_frame_line_pixel_5_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_5_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_5_2[7:0]  ), //i
    .ab       (sIMD2INT8_1157_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1157_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1158 (
    .a        (prevConv_payload_frame_line_pixel_6_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_6_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_6_2[7:0]  ), //i
    .ab       (sIMD2INT8_1158_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1158_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1159 (
    .a        (prevConv_payload_frame_line_pixel_7_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_7_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_7_2[7:0]  ), //i
    .ab       (sIMD2INT8_1159_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1159_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1160 (
    .a        (prevConv_payload_frame_line_pixel_8_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_8_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_8_2[7:0]  ), //i
    .ab       (sIMD2INT8_1160_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1160_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1161 (
    .a        (prevConv_payload_frame_line_pixel_9_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_9_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_9_2[7:0]  ), //i
    .ab       (sIMD2INT8_1161_ab[15:0]                     ), //o
    .ac       (sIMD2INT8_1161_ac[15:0]                     ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                       ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                       ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                       ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                       ), //i
    .clk      (clk                                         )  //i
  );
  SIMD2INT8 sIMD2INT8_1162 (
    .a        (prevConv_payload_frame_line_pixel_10_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_10_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_10_2[7:0]  ), //i
    .ab       (sIMD2INT8_1162_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1162_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1163 (
    .a        (prevConv_payload_frame_line_pixel_11_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_11_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_11_2[7:0]  ), //i
    .ab       (sIMD2INT8_1163_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1163_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1164 (
    .a        (prevConv_payload_frame_line_pixel_12_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_12_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_12_2[7:0]  ), //i
    .ab       (sIMD2INT8_1164_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1164_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1165 (
    .a        (prevConv_payload_frame_line_pixel_13_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_13_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_13_2[7:0]  ), //i
    .ab       (sIMD2INT8_1165_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1165_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1166 (
    .a        (prevConv_payload_frame_line_pixel_14_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_14_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_14_2[7:0]  ), //i
    .ab       (sIMD2INT8_1166_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1166_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1167 (
    .a        (prevConv_payload_frame_line_pixel_15_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_15_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_15_2[7:0]  ), //i
    .ab       (sIMD2INT8_1167_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1167_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1168 (
    .a        (prevConv_payload_frame_line_pixel_16_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_16_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_16_2[7:0]  ), //i
    .ab       (sIMD2INT8_1168_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1168_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1169 (
    .a        (prevConv_payload_frame_line_pixel_17_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_17_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_17_2[7:0]  ), //i
    .ab       (sIMD2INT8_1169_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1169_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1170 (
    .a        (prevConv_payload_frame_line_pixel_18_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_18_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_18_2[7:0]  ), //i
    .ab       (sIMD2INT8_1170_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1170_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1171 (
    .a        (prevConv_payload_frame_line_pixel_19_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_19_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_19_2[7:0]  ), //i
    .ab       (sIMD2INT8_1171_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1171_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1172 (
    .a        (prevConv_payload_frame_line_pixel_20_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_20_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_20_2[7:0]  ), //i
    .ab       (sIMD2INT8_1172_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1172_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1173 (
    .a        (prevConv_payload_frame_line_pixel_21_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_21_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_21_2[7:0]  ), //i
    .ab       (sIMD2INT8_1173_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1173_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1174 (
    .a        (prevConv_payload_frame_line_pixel_22_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_22_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_22_2[7:0]  ), //i
    .ab       (sIMD2INT8_1174_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1174_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1175 (
    .a        (prevConv_payload_frame_line_pixel_23_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_23_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_23_2[7:0]  ), //i
    .ab       (sIMD2INT8_1175_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1175_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1176 (
    .a        (prevConv_payload_frame_line_pixel_24_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_24_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_24_2[7:0]  ), //i
    .ab       (sIMD2INT8_1176_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1176_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1177 (
    .a        (prevConv_payload_frame_line_pixel_25_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_25_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_25_2[7:0]  ), //i
    .ab       (sIMD2INT8_1177_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1177_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1178 (
    .a        (prevConv_payload_frame_line_pixel_26_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_26_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_26_2[7:0]  ), //i
    .ab       (sIMD2INT8_1178_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1178_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1179 (
    .a        (prevConv_payload_frame_line_pixel_27_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_27_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_27_2[7:0]  ), //i
    .ab       (sIMD2INT8_1179_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1179_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1180 (
    .a        (prevConv_payload_frame_line_pixel_28_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_28_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_28_2[7:0]  ), //i
    .ab       (sIMD2INT8_1180_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1180_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1181 (
    .a        (prevConv_payload_frame_line_pixel_29_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_29_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_29_2[7:0]  ), //i
    .ab       (sIMD2INT8_1181_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1181_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1182 (
    .a        (prevConv_payload_frame_line_pixel_30_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_30_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_30_2[7:0]  ), //i
    .ab       (sIMD2INT8_1182_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1182_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1183 (
    .a        (prevConv_payload_frame_line_pixel_31_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_31_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_31_2[7:0]  ), //i
    .ab       (sIMD2INT8_1183_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1183_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1184 (
    .a        (prevConv_payload_frame_line_pixel_32_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_32_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_32_2[7:0]  ), //i
    .ab       (sIMD2INT8_1184_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1184_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1185 (
    .a        (prevConv_payload_frame_line_pixel_33_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_33_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_33_2[7:0]  ), //i
    .ab       (sIMD2INT8_1185_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1185_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1186 (
    .a        (prevConv_payload_frame_line_pixel_34_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_34_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_34_2[7:0]  ), //i
    .ab       (sIMD2INT8_1186_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1186_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1187 (
    .a        (prevConv_payload_frame_line_pixel_35_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_35_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_35_2[7:0]  ), //i
    .ab       (sIMD2INT8_1187_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1187_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1188 (
    .a        (prevConv_payload_frame_line_pixel_36_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_36_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_36_2[7:0]  ), //i
    .ab       (sIMD2INT8_1188_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1188_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1189 (
    .a        (prevConv_payload_frame_line_pixel_37_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_37_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_37_2[7:0]  ), //i
    .ab       (sIMD2INT8_1189_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1189_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1190 (
    .a        (prevConv_payload_frame_line_pixel_38_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_38_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_38_2[7:0]  ), //i
    .ab       (sIMD2INT8_1190_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1190_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1191 (
    .a        (prevConv_payload_frame_line_pixel_39_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_39_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_39_2[7:0]  ), //i
    .ab       (sIMD2INT8_1191_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1191_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1192 (
    .a        (prevConv_payload_frame_line_pixel_40_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_40_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_40_2[7:0]  ), //i
    .ab       (sIMD2INT8_1192_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1192_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1193 (
    .a        (prevConv_payload_frame_line_pixel_41_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_41_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_41_2[7:0]  ), //i
    .ab       (sIMD2INT8_1193_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1193_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1194 (
    .a        (prevConv_payload_frame_line_pixel_42_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_42_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_42_2[7:0]  ), //i
    .ab       (sIMD2INT8_1194_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1194_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1195 (
    .a        (prevConv_payload_frame_line_pixel_43_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_43_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_43_2[7:0]  ), //i
    .ab       (sIMD2INT8_1195_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1195_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1196 (
    .a        (prevConv_payload_frame_line_pixel_44_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_44_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_44_2[7:0]  ), //i
    .ab       (sIMD2INT8_1196_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1196_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1197 (
    .a        (prevConv_payload_frame_line_pixel_45_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_45_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_45_2[7:0]  ), //i
    .ab       (sIMD2INT8_1197_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1197_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1198 (
    .a        (prevConv_payload_frame_line_pixel_46_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_46_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_46_2[7:0]  ), //i
    .ab       (sIMD2INT8_1198_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1198_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1199 (
    .a        (prevConv_payload_frame_line_pixel_47_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_47_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_47_2[7:0]  ), //i
    .ab       (sIMD2INT8_1199_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1199_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1200 (
    .a        (prevConv_payload_frame_line_pixel_48_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_48_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_48_2[7:0]  ), //i
    .ab       (sIMD2INT8_1200_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1200_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1201 (
    .a        (prevConv_payload_frame_line_pixel_49_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_49_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_49_2[7:0]  ), //i
    .ab       (sIMD2INT8_1201_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1201_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1202 (
    .a        (prevConv_payload_frame_line_pixel_50_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_50_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_50_2[7:0]  ), //i
    .ab       (sIMD2INT8_1202_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1202_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1203 (
    .a        (prevConv_payload_frame_line_pixel_51_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_51_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_51_2[7:0]  ), //i
    .ab       (sIMD2INT8_1203_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1203_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1204 (
    .a        (prevConv_payload_frame_line_pixel_52_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_52_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_52_2[7:0]  ), //i
    .ab       (sIMD2INT8_1204_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1204_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1205 (
    .a        (prevConv_payload_frame_line_pixel_53_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_53_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_53_2[7:0]  ), //i
    .ab       (sIMD2INT8_1205_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1205_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1206 (
    .a        (prevConv_payload_frame_line_pixel_54_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_54_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_54_2[7:0]  ), //i
    .ab       (sIMD2INT8_1206_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1206_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1207 (
    .a        (prevConv_payload_frame_line_pixel_55_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_55_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_55_2[7:0]  ), //i
    .ab       (sIMD2INT8_1207_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1207_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1208 (
    .a        (prevConv_payload_frame_line_pixel_56_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_56_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_56_2[7:0]  ), //i
    .ab       (sIMD2INT8_1208_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1208_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1209 (
    .a        (prevConv_payload_frame_line_pixel_57_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_57_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_57_2[7:0]  ), //i
    .ab       (sIMD2INT8_1209_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1209_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1210 (
    .a        (prevConv_payload_frame_line_pixel_58_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_58_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_58_2[7:0]  ), //i
    .ab       (sIMD2INT8_1210_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1210_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1211 (
    .a        (prevConv_payload_frame_line_pixel_59_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_59_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_59_2[7:0]  ), //i
    .ab       (sIMD2INT8_1211_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1211_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1212 (
    .a        (prevConv_payload_frame_line_pixel_60_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_60_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_60_2[7:0]  ), //i
    .ab       (sIMD2INT8_1212_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1212_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1213 (
    .a        (prevConv_payload_frame_line_pixel_61_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_61_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_61_2[7:0]  ), //i
    .ab       (sIMD2INT8_1213_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1213_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1214 (
    .a        (prevConv_payload_frame_line_pixel_62_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_62_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_62_2[7:0]  ), //i
    .ab       (sIMD2INT8_1214_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1214_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1215 (
    .a        (prevConv_payload_frame_line_pixel_63_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_63_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_63_2[7:0]  ), //i
    .ab       (sIMD2INT8_1215_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1215_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1216 (
    .a        (prevConv_payload_frame_line_pixel_64_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_64_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_64_2[7:0]  ), //i
    .ab       (sIMD2INT8_1216_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1216_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1217 (
    .a        (prevConv_payload_frame_line_pixel_65_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_65_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_65_2[7:0]  ), //i
    .ab       (sIMD2INT8_1217_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1217_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1218 (
    .a        (prevConv_payload_frame_line_pixel_66_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_66_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_66_2[7:0]  ), //i
    .ab       (sIMD2INT8_1218_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1218_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1219 (
    .a        (prevConv_payload_frame_line_pixel_67_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_67_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_67_2[7:0]  ), //i
    .ab       (sIMD2INT8_1219_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1219_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1220 (
    .a        (prevConv_payload_frame_line_pixel_68_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_68_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_68_2[7:0]  ), //i
    .ab       (sIMD2INT8_1220_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1220_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1221 (
    .a        (prevConv_payload_frame_line_pixel_69_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_69_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_69_2[7:0]  ), //i
    .ab       (sIMD2INT8_1221_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1221_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1222 (
    .a        (prevConv_payload_frame_line_pixel_70_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_70_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_70_2[7:0]  ), //i
    .ab       (sIMD2INT8_1222_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1222_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1223 (
    .a        (prevConv_payload_frame_line_pixel_71_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_71_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_71_2[7:0]  ), //i
    .ab       (sIMD2INT8_1223_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1223_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1224 (
    .a        (prevConv_payload_frame_line_pixel_72_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_72_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_72_2[7:0]  ), //i
    .ab       (sIMD2INT8_1224_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1224_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1225 (
    .a        (prevConv_payload_frame_line_pixel_73_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_73_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_73_2[7:0]  ), //i
    .ab       (sIMD2INT8_1225_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1225_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1226 (
    .a        (prevConv_payload_frame_line_pixel_74_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_74_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_74_2[7:0]  ), //i
    .ab       (sIMD2INT8_1226_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1226_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1227 (
    .a        (prevConv_payload_frame_line_pixel_75_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_75_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_75_2[7:0]  ), //i
    .ab       (sIMD2INT8_1227_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1227_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1228 (
    .a        (prevConv_payload_frame_line_pixel_76_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_76_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_76_2[7:0]  ), //i
    .ab       (sIMD2INT8_1228_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1228_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1229 (
    .a        (prevConv_payload_frame_line_pixel_77_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_77_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_77_2[7:0]  ), //i
    .ab       (sIMD2INT8_1229_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1229_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1230 (
    .a        (prevConv_payload_frame_line_pixel_78_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_78_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_78_2[7:0]  ), //i
    .ab       (sIMD2INT8_1230_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1230_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1231 (
    .a        (prevConv_payload_frame_line_pixel_79_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_79_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_79_2[7:0]  ), //i
    .ab       (sIMD2INT8_1231_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1231_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1232 (
    .a        (prevConv_payload_frame_line_pixel_80_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_80_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_80_2[7:0]  ), //i
    .ab       (sIMD2INT8_1232_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1232_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1233 (
    .a        (prevConv_payload_frame_line_pixel_81_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_81_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_81_2[7:0]  ), //i
    .ab       (sIMD2INT8_1233_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1233_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1234 (
    .a        (prevConv_payload_frame_line_pixel_82_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_82_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_82_2[7:0]  ), //i
    .ab       (sIMD2INT8_1234_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1234_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1235 (
    .a        (prevConv_payload_frame_line_pixel_83_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_83_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_83_2[7:0]  ), //i
    .ab       (sIMD2INT8_1235_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1235_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1236 (
    .a        (prevConv_payload_frame_line_pixel_84_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_84_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_84_2[7:0]  ), //i
    .ab       (sIMD2INT8_1236_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1236_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1237 (
    .a        (prevConv_payload_frame_line_pixel_85_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_85_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_85_2[7:0]  ), //i
    .ab       (sIMD2INT8_1237_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1237_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1238 (
    .a        (prevConv_payload_frame_line_pixel_86_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_86_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_86_2[7:0]  ), //i
    .ab       (sIMD2INT8_1238_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1238_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1239 (
    .a        (prevConv_payload_frame_line_pixel_87_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_87_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_87_2[7:0]  ), //i
    .ab       (sIMD2INT8_1239_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1239_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1240 (
    .a        (prevConv_payload_frame_line_pixel_88_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_88_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_88_2[7:0]  ), //i
    .ab       (sIMD2INT8_1240_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1240_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1241 (
    .a        (prevConv_payload_frame_line_pixel_89_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_89_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_89_2[7:0]  ), //i
    .ab       (sIMD2INT8_1241_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1241_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1242 (
    .a        (prevConv_payload_frame_line_pixel_90_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_90_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_90_2[7:0]  ), //i
    .ab       (sIMD2INT8_1242_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1242_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1243 (
    .a        (prevConv_payload_frame_line_pixel_91_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_91_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_91_2[7:0]  ), //i
    .ab       (sIMD2INT8_1243_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1243_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1244 (
    .a        (prevConv_payload_frame_line_pixel_92_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_92_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_92_2[7:0]  ), //i
    .ab       (sIMD2INT8_1244_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1244_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1245 (
    .a        (prevConv_payload_frame_line_pixel_93_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_93_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_93_2[7:0]  ), //i
    .ab       (sIMD2INT8_1245_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1245_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1246 (
    .a        (prevConv_payload_frame_line_pixel_94_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_94_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_94_2[7:0]  ), //i
    .ab       (sIMD2INT8_1246_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1246_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1247 (
    .a        (prevConv_payload_frame_line_pixel_95_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_95_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_95_2[7:0]  ), //i
    .ab       (sIMD2INT8_1247_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1247_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1248 (
    .a        (prevConv_payload_frame_line_pixel_96_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_96_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_96_2[7:0]  ), //i
    .ab       (sIMD2INT8_1248_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1248_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1249 (
    .a        (prevConv_payload_frame_line_pixel_97_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_97_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_97_2[7:0]  ), //i
    .ab       (sIMD2INT8_1249_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1249_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1250 (
    .a        (prevConv_payload_frame_line_pixel_98_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_98_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_98_2[7:0]  ), //i
    .ab       (sIMD2INT8_1250_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1250_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1251 (
    .a        (prevConv_payload_frame_line_pixel_99_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_99_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_99_2[7:0]  ), //i
    .ab       (sIMD2INT8_1251_ab[15:0]                      ), //o
    .ac       (sIMD2INT8_1251_ac[15:0]                      ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                        ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                        ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                        ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                        ), //i
    .clk      (clk                                          )  //i
  );
  SIMD2INT8 sIMD2INT8_1252 (
    .a        (prevConv_payload_frame_line_pixel_100_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_100_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_100_2[7:0]  ), //i
    .ab       (sIMD2INT8_1252_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1252_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1253 (
    .a        (prevConv_payload_frame_line_pixel_101_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_101_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_101_2[7:0]  ), //i
    .ab       (sIMD2INT8_1253_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1253_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1254 (
    .a        (prevConv_payload_frame_line_pixel_102_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_102_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_102_2[7:0]  ), //i
    .ab       (sIMD2INT8_1254_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1254_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1255 (
    .a        (prevConv_payload_frame_line_pixel_103_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_103_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_103_2[7:0]  ), //i
    .ab       (sIMD2INT8_1255_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1255_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1256 (
    .a        (prevConv_payload_frame_line_pixel_104_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_104_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_104_2[7:0]  ), //i
    .ab       (sIMD2INT8_1256_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1256_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1257 (
    .a        (prevConv_payload_frame_line_pixel_105_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_105_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_105_2[7:0]  ), //i
    .ab       (sIMD2INT8_1257_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1257_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1258 (
    .a        (prevConv_payload_frame_line_pixel_106_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_106_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_106_2[7:0]  ), //i
    .ab       (sIMD2INT8_1258_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1258_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1259 (
    .a        (prevConv_payload_frame_line_pixel_107_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_107_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_107_2[7:0]  ), //i
    .ab       (sIMD2INT8_1259_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1259_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1260 (
    .a        (prevConv_payload_frame_line_pixel_108_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_108_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_108_2[7:0]  ), //i
    .ab       (sIMD2INT8_1260_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1260_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1261 (
    .a        (prevConv_payload_frame_line_pixel_109_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_109_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_109_2[7:0]  ), //i
    .ab       (sIMD2INT8_1261_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1261_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1262 (
    .a        (prevConv_payload_frame_line_pixel_110_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_110_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_110_2[7:0]  ), //i
    .ab       (sIMD2INT8_1262_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1262_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1263 (
    .a        (prevConv_payload_frame_line_pixel_111_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_111_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_111_2[7:0]  ), //i
    .ab       (sIMD2INT8_1263_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1263_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1264 (
    .a        (prevConv_payload_frame_line_pixel_112_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_112_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_112_2[7:0]  ), //i
    .ab       (sIMD2INT8_1264_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1264_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1265 (
    .a        (prevConv_payload_frame_line_pixel_113_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_113_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_113_2[7:0]  ), //i
    .ab       (sIMD2INT8_1265_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1265_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1266 (
    .a        (prevConv_payload_frame_line_pixel_114_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_114_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_114_2[7:0]  ), //i
    .ab       (sIMD2INT8_1266_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1266_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1267 (
    .a        (prevConv_payload_frame_line_pixel_115_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_115_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_115_2[7:0]  ), //i
    .ab       (sIMD2INT8_1267_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1267_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1268 (
    .a        (prevConv_payload_frame_line_pixel_116_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_116_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_116_2[7:0]  ), //i
    .ab       (sIMD2INT8_1268_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1268_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1269 (
    .a        (prevConv_payload_frame_line_pixel_117_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_117_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_117_2[7:0]  ), //i
    .ab       (sIMD2INT8_1269_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1269_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1270 (
    .a        (prevConv_payload_frame_line_pixel_118_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_118_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_118_2[7:0]  ), //i
    .ab       (sIMD2INT8_1270_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1270_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1271 (
    .a        (prevConv_payload_frame_line_pixel_119_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_119_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_119_2[7:0]  ), //i
    .ab       (sIMD2INT8_1271_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1271_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1272 (
    .a        (prevConv_payload_frame_line_pixel_120_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_120_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_120_2[7:0]  ), //i
    .ab       (sIMD2INT8_1272_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1272_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1273 (
    .a        (prevConv_payload_frame_line_pixel_121_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_121_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_121_2[7:0]  ), //i
    .ab       (sIMD2INT8_1273_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1273_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1274 (
    .a        (prevConv_payload_frame_line_pixel_122_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_122_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_122_2[7:0]  ), //i
    .ab       (sIMD2INT8_1274_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1274_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1275 (
    .a        (prevConv_payload_frame_line_pixel_123_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_123_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_123_2[7:0]  ), //i
    .ab       (sIMD2INT8_1275_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1275_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1276 (
    .a        (prevConv_payload_frame_line_pixel_124_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_124_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_124_2[7:0]  ), //i
    .ab       (sIMD2INT8_1276_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1276_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1277 (
    .a        (prevConv_payload_frame_line_pixel_125_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_125_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_125_2[7:0]  ), //i
    .ab       (sIMD2INT8_1277_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1277_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1278 (
    .a        (prevConv_payload_frame_line_pixel_126_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_126_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_126_2[7:0]  ), //i
    .ab       (sIMD2INT8_1278_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1278_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1279 (
    .a        (prevConv_payload_frame_line_pixel_127_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_127_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_127_2[7:0]  ), //i
    .ab       (sIMD2INT8_1279_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1279_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1280 (
    .a        (prevConv_payload_frame_line_pixel_128_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_128_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_128_2[7:0]  ), //i
    .ab       (sIMD2INT8_1280_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1280_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1281 (
    .a        (prevConv_payload_frame_line_pixel_129_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_129_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_129_2[7:0]  ), //i
    .ab       (sIMD2INT8_1281_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1281_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1282 (
    .a        (prevConv_payload_frame_line_pixel_130_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_130_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_130_2[7:0]  ), //i
    .ab       (sIMD2INT8_1282_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1282_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1283 (
    .a        (prevConv_payload_frame_line_pixel_131_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_131_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_131_2[7:0]  ), //i
    .ab       (sIMD2INT8_1283_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1283_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1284 (
    .a        (prevConv_payload_frame_line_pixel_132_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_132_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_132_2[7:0]  ), //i
    .ab       (sIMD2INT8_1284_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1284_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1285 (
    .a        (prevConv_payload_frame_line_pixel_133_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_133_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_133_2[7:0]  ), //i
    .ab       (sIMD2INT8_1285_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1285_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1286 (
    .a        (prevConv_payload_frame_line_pixel_134_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_134_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_134_2[7:0]  ), //i
    .ab       (sIMD2INT8_1286_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1286_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1287 (
    .a        (prevConv_payload_frame_line_pixel_135_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_135_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_135_2[7:0]  ), //i
    .ab       (sIMD2INT8_1287_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1287_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1288 (
    .a        (prevConv_payload_frame_line_pixel_136_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_136_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_136_2[7:0]  ), //i
    .ab       (sIMD2INT8_1288_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1288_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1289 (
    .a        (prevConv_payload_frame_line_pixel_137_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_137_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_137_2[7:0]  ), //i
    .ab       (sIMD2INT8_1289_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1289_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1290 (
    .a        (prevConv_payload_frame_line_pixel_138_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_138_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_138_2[7:0]  ), //i
    .ab       (sIMD2INT8_1290_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1290_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1291 (
    .a        (prevConv_payload_frame_line_pixel_139_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_139_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_139_2[7:0]  ), //i
    .ab       (sIMD2INT8_1291_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1291_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1292 (
    .a        (prevConv_payload_frame_line_pixel_140_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_140_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_140_2[7:0]  ), //i
    .ab       (sIMD2INT8_1292_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1292_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1293 (
    .a        (prevConv_payload_frame_line_pixel_141_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_141_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_141_2[7:0]  ), //i
    .ab       (sIMD2INT8_1293_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1293_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1294 (
    .a        (prevConv_payload_frame_line_pixel_142_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_142_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_142_2[7:0]  ), //i
    .ab       (sIMD2INT8_1294_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1294_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  SIMD2INT8 sIMD2INT8_1295 (
    .a        (prevConv_payload_frame_line_pixel_143_0[7:0]  ), //i
    .b        (prevConv_payload_frame_line_pixel_143_1[7:0]  ), //i
    .c        (prevConv_payload_frame_line_pixel_143_2[7:0]  ), //i
    .ab       (sIMD2INT8_1295_ab[15:0]                       ), //o
    .ac       (sIMD2INT8_1295_ac[15:0]                       ), //o
    .CEs_0    (eventM2sPipes_9_CEs_0                         ), //i
    .CEs_1    (eventM2sPipes_9_CEs_1                         ), //i
    .CEs_2    (eventM2sPipes_9_CEs_2                         ), //i
    .CEs_3    (eventM2sPipes_9_CEs_3                         ), //i
    .clk      (clk                                           )  //i
  );
  VideoFrameHistory acc (
    .numberOfInputFrames                      (numberOfInputFrames[7:0]                           ), //i
    .numberOfOutputFrames                     (numberOfOutputFrames[7:0]                          ), //i
    .videoIn_valid                            (postConv_s2mPipe_valid                             ), //i
    .videoIn_ready                            (acc_videoIn_ready                                  ), //o
    .videoIn_payload_frame_line_pixel_0       (postConv_s2mPipe_payload_frame_line_pixel_0[15:0]  ), //i
    .videoIn_payload_frame_line_pixel_1       (postConv_s2mPipe_payload_frame_line_pixel_1[15:0]  ), //i
    .videoIn_payload_frame_line_endOfLine     (postConv_s2mPipe_payload_frame_line_endOfLine      ), //i
    .videoIn_payload_frame_endOfFrame         (postConv_s2mPipe_payload_frame_endOfFrame          ), //i
    .videoIn_payload_endOfPack                (postConv_s2mPipe_payload_endOfPack                 ), //i
    .videoOut_valid                           (acc_videoOut_valid                                 ), //o
    .videoOut_ready                           (outputs_ready                                      ), //i
    .videoOut_payload_frame_line_pixel_0      (acc_videoOut_payload_frame_line_pixel_0[23:0]      ), //o
    .videoOut_payload_frame_line_pixel_1      (acc_videoOut_payload_frame_line_pixel_1[23:0]      ), //o
    .videoOut_payload_frame_line_endOfLine    (acc_videoOut_payload_frame_line_endOfLine          ), //o
    .videoOut_payload_frame_endOfFrame        (acc_videoOut_payload_frame_endOfFrame              ), //o
    .videoOut_payload_endOfPack               (acc_videoOut_payload_endOfPack                     ), //o
    .clk                                      (clk                                                ), //i
    .reset                                    (reset                                              )  //i
  );
  assign tmp_inputs_ready = (! (! weights_valid));
  assign inputsT_valid = (inputs_valid && tmp_inputs_ready);
  assign inputs_ready = (inputsT_ready && tmp_inputs_ready);
  assign inputsT_payload_frame_line_pixel_0_0_0 = inputs_payload_frame_line_pixel_0_0_0;
  assign inputsT_payload_frame_line_pixel_0_0_1 = inputs_payload_frame_line_pixel_0_0_1;
  assign inputsT_payload_frame_line_pixel_0_0_2 = inputs_payload_frame_line_pixel_0_0_2;
  assign inputsT_payload_frame_line_pixel_0_0_3 = inputs_payload_frame_line_pixel_0_0_3;
  assign inputsT_payload_frame_line_pixel_0_0_4 = inputs_payload_frame_line_pixel_0_0_4;
  assign inputsT_payload_frame_line_pixel_0_0_5 = inputs_payload_frame_line_pixel_0_0_5;
  assign inputsT_payload_frame_line_pixel_0_0_6 = inputs_payload_frame_line_pixel_0_0_6;
  assign inputsT_payload_frame_line_pixel_0_0_7 = inputs_payload_frame_line_pixel_0_0_7;
  assign inputsT_payload_frame_line_pixel_0_0_8 = inputs_payload_frame_line_pixel_0_0_8;
  assign inputsT_payload_frame_line_pixel_0_0_9 = inputs_payload_frame_line_pixel_0_0_9;
  assign inputsT_payload_frame_line_pixel_0_0_10 = inputs_payload_frame_line_pixel_0_0_10;
  assign inputsT_payload_frame_line_pixel_0_0_11 = inputs_payload_frame_line_pixel_0_0_11;
  assign inputsT_payload_frame_line_pixel_0_0_12 = inputs_payload_frame_line_pixel_0_0_12;
  assign inputsT_payload_frame_line_pixel_0_0_13 = inputs_payload_frame_line_pixel_0_0_13;
  assign inputsT_payload_frame_line_pixel_0_0_14 = inputs_payload_frame_line_pixel_0_0_14;
  assign inputsT_payload_frame_line_pixel_0_0_15 = inputs_payload_frame_line_pixel_0_0_15;
  assign inputsT_payload_frame_line_pixel_0_1_0 = inputs_payload_frame_line_pixel_0_1_0;
  assign inputsT_payload_frame_line_pixel_0_1_1 = inputs_payload_frame_line_pixel_0_1_1;
  assign inputsT_payload_frame_line_pixel_0_1_2 = inputs_payload_frame_line_pixel_0_1_2;
  assign inputsT_payload_frame_line_pixel_0_1_3 = inputs_payload_frame_line_pixel_0_1_3;
  assign inputsT_payload_frame_line_pixel_0_1_4 = inputs_payload_frame_line_pixel_0_1_4;
  assign inputsT_payload_frame_line_pixel_0_1_5 = inputs_payload_frame_line_pixel_0_1_5;
  assign inputsT_payload_frame_line_pixel_0_1_6 = inputs_payload_frame_line_pixel_0_1_6;
  assign inputsT_payload_frame_line_pixel_0_1_7 = inputs_payload_frame_line_pixel_0_1_7;
  assign inputsT_payload_frame_line_pixel_0_1_8 = inputs_payload_frame_line_pixel_0_1_8;
  assign inputsT_payload_frame_line_pixel_0_1_9 = inputs_payload_frame_line_pixel_0_1_9;
  assign inputsT_payload_frame_line_pixel_0_1_10 = inputs_payload_frame_line_pixel_0_1_10;
  assign inputsT_payload_frame_line_pixel_0_1_11 = inputs_payload_frame_line_pixel_0_1_11;
  assign inputsT_payload_frame_line_pixel_0_1_12 = inputs_payload_frame_line_pixel_0_1_12;
  assign inputsT_payload_frame_line_pixel_0_1_13 = inputs_payload_frame_line_pixel_0_1_13;
  assign inputsT_payload_frame_line_pixel_0_1_14 = inputs_payload_frame_line_pixel_0_1_14;
  assign inputsT_payload_frame_line_pixel_0_1_15 = inputs_payload_frame_line_pixel_0_1_15;
  assign inputsT_payload_frame_line_pixel_0_2_0 = inputs_payload_frame_line_pixel_0_2_0;
  assign inputsT_payload_frame_line_pixel_0_2_1 = inputs_payload_frame_line_pixel_0_2_1;
  assign inputsT_payload_frame_line_pixel_0_2_2 = inputs_payload_frame_line_pixel_0_2_2;
  assign inputsT_payload_frame_line_pixel_0_2_3 = inputs_payload_frame_line_pixel_0_2_3;
  assign inputsT_payload_frame_line_pixel_0_2_4 = inputs_payload_frame_line_pixel_0_2_4;
  assign inputsT_payload_frame_line_pixel_0_2_5 = inputs_payload_frame_line_pixel_0_2_5;
  assign inputsT_payload_frame_line_pixel_0_2_6 = inputs_payload_frame_line_pixel_0_2_6;
  assign inputsT_payload_frame_line_pixel_0_2_7 = inputs_payload_frame_line_pixel_0_2_7;
  assign inputsT_payload_frame_line_pixel_0_2_8 = inputs_payload_frame_line_pixel_0_2_8;
  assign inputsT_payload_frame_line_pixel_0_2_9 = inputs_payload_frame_line_pixel_0_2_9;
  assign inputsT_payload_frame_line_pixel_0_2_10 = inputs_payload_frame_line_pixel_0_2_10;
  assign inputsT_payload_frame_line_pixel_0_2_11 = inputs_payload_frame_line_pixel_0_2_11;
  assign inputsT_payload_frame_line_pixel_0_2_12 = inputs_payload_frame_line_pixel_0_2_12;
  assign inputsT_payload_frame_line_pixel_0_2_13 = inputs_payload_frame_line_pixel_0_2_13;
  assign inputsT_payload_frame_line_pixel_0_2_14 = inputs_payload_frame_line_pixel_0_2_14;
  assign inputsT_payload_frame_line_pixel_0_2_15 = inputs_payload_frame_line_pixel_0_2_15;
  assign inputsT_payload_frame_line_pixel_1_0_0 = inputs_payload_frame_line_pixel_1_0_0;
  assign inputsT_payload_frame_line_pixel_1_0_1 = inputs_payload_frame_line_pixel_1_0_1;
  assign inputsT_payload_frame_line_pixel_1_0_2 = inputs_payload_frame_line_pixel_1_0_2;
  assign inputsT_payload_frame_line_pixel_1_0_3 = inputs_payload_frame_line_pixel_1_0_3;
  assign inputsT_payload_frame_line_pixel_1_0_4 = inputs_payload_frame_line_pixel_1_0_4;
  assign inputsT_payload_frame_line_pixel_1_0_5 = inputs_payload_frame_line_pixel_1_0_5;
  assign inputsT_payload_frame_line_pixel_1_0_6 = inputs_payload_frame_line_pixel_1_0_6;
  assign inputsT_payload_frame_line_pixel_1_0_7 = inputs_payload_frame_line_pixel_1_0_7;
  assign inputsT_payload_frame_line_pixel_1_0_8 = inputs_payload_frame_line_pixel_1_0_8;
  assign inputsT_payload_frame_line_pixel_1_0_9 = inputs_payload_frame_line_pixel_1_0_9;
  assign inputsT_payload_frame_line_pixel_1_0_10 = inputs_payload_frame_line_pixel_1_0_10;
  assign inputsT_payload_frame_line_pixel_1_0_11 = inputs_payload_frame_line_pixel_1_0_11;
  assign inputsT_payload_frame_line_pixel_1_0_12 = inputs_payload_frame_line_pixel_1_0_12;
  assign inputsT_payload_frame_line_pixel_1_0_13 = inputs_payload_frame_line_pixel_1_0_13;
  assign inputsT_payload_frame_line_pixel_1_0_14 = inputs_payload_frame_line_pixel_1_0_14;
  assign inputsT_payload_frame_line_pixel_1_0_15 = inputs_payload_frame_line_pixel_1_0_15;
  assign inputsT_payload_frame_line_pixel_1_1_0 = inputs_payload_frame_line_pixel_1_1_0;
  assign inputsT_payload_frame_line_pixel_1_1_1 = inputs_payload_frame_line_pixel_1_1_1;
  assign inputsT_payload_frame_line_pixel_1_1_2 = inputs_payload_frame_line_pixel_1_1_2;
  assign inputsT_payload_frame_line_pixel_1_1_3 = inputs_payload_frame_line_pixel_1_1_3;
  assign inputsT_payload_frame_line_pixel_1_1_4 = inputs_payload_frame_line_pixel_1_1_4;
  assign inputsT_payload_frame_line_pixel_1_1_5 = inputs_payload_frame_line_pixel_1_1_5;
  assign inputsT_payload_frame_line_pixel_1_1_6 = inputs_payload_frame_line_pixel_1_1_6;
  assign inputsT_payload_frame_line_pixel_1_1_7 = inputs_payload_frame_line_pixel_1_1_7;
  assign inputsT_payload_frame_line_pixel_1_1_8 = inputs_payload_frame_line_pixel_1_1_8;
  assign inputsT_payload_frame_line_pixel_1_1_9 = inputs_payload_frame_line_pixel_1_1_9;
  assign inputsT_payload_frame_line_pixel_1_1_10 = inputs_payload_frame_line_pixel_1_1_10;
  assign inputsT_payload_frame_line_pixel_1_1_11 = inputs_payload_frame_line_pixel_1_1_11;
  assign inputsT_payload_frame_line_pixel_1_1_12 = inputs_payload_frame_line_pixel_1_1_12;
  assign inputsT_payload_frame_line_pixel_1_1_13 = inputs_payload_frame_line_pixel_1_1_13;
  assign inputsT_payload_frame_line_pixel_1_1_14 = inputs_payload_frame_line_pixel_1_1_14;
  assign inputsT_payload_frame_line_pixel_1_1_15 = inputs_payload_frame_line_pixel_1_1_15;
  assign inputsT_payload_frame_line_pixel_1_2_0 = inputs_payload_frame_line_pixel_1_2_0;
  assign inputsT_payload_frame_line_pixel_1_2_1 = inputs_payload_frame_line_pixel_1_2_1;
  assign inputsT_payload_frame_line_pixel_1_2_2 = inputs_payload_frame_line_pixel_1_2_2;
  assign inputsT_payload_frame_line_pixel_1_2_3 = inputs_payload_frame_line_pixel_1_2_3;
  assign inputsT_payload_frame_line_pixel_1_2_4 = inputs_payload_frame_line_pixel_1_2_4;
  assign inputsT_payload_frame_line_pixel_1_2_5 = inputs_payload_frame_line_pixel_1_2_5;
  assign inputsT_payload_frame_line_pixel_1_2_6 = inputs_payload_frame_line_pixel_1_2_6;
  assign inputsT_payload_frame_line_pixel_1_2_7 = inputs_payload_frame_line_pixel_1_2_7;
  assign inputsT_payload_frame_line_pixel_1_2_8 = inputs_payload_frame_line_pixel_1_2_8;
  assign inputsT_payload_frame_line_pixel_1_2_9 = inputs_payload_frame_line_pixel_1_2_9;
  assign inputsT_payload_frame_line_pixel_1_2_10 = inputs_payload_frame_line_pixel_1_2_10;
  assign inputsT_payload_frame_line_pixel_1_2_11 = inputs_payload_frame_line_pixel_1_2_11;
  assign inputsT_payload_frame_line_pixel_1_2_12 = inputs_payload_frame_line_pixel_1_2_12;
  assign inputsT_payload_frame_line_pixel_1_2_13 = inputs_payload_frame_line_pixel_1_2_13;
  assign inputsT_payload_frame_line_pixel_1_2_14 = inputs_payload_frame_line_pixel_1_2_14;
  assign inputsT_payload_frame_line_pixel_1_2_15 = inputs_payload_frame_line_pixel_1_2_15;
  assign inputsT_payload_frame_line_pixel_2_0_0 = inputs_payload_frame_line_pixel_2_0_0;
  assign inputsT_payload_frame_line_pixel_2_0_1 = inputs_payload_frame_line_pixel_2_0_1;
  assign inputsT_payload_frame_line_pixel_2_0_2 = inputs_payload_frame_line_pixel_2_0_2;
  assign inputsT_payload_frame_line_pixel_2_0_3 = inputs_payload_frame_line_pixel_2_0_3;
  assign inputsT_payload_frame_line_pixel_2_0_4 = inputs_payload_frame_line_pixel_2_0_4;
  assign inputsT_payload_frame_line_pixel_2_0_5 = inputs_payload_frame_line_pixel_2_0_5;
  assign inputsT_payload_frame_line_pixel_2_0_6 = inputs_payload_frame_line_pixel_2_0_6;
  assign inputsT_payload_frame_line_pixel_2_0_7 = inputs_payload_frame_line_pixel_2_0_7;
  assign inputsT_payload_frame_line_pixel_2_0_8 = inputs_payload_frame_line_pixel_2_0_8;
  assign inputsT_payload_frame_line_pixel_2_0_9 = inputs_payload_frame_line_pixel_2_0_9;
  assign inputsT_payload_frame_line_pixel_2_0_10 = inputs_payload_frame_line_pixel_2_0_10;
  assign inputsT_payload_frame_line_pixel_2_0_11 = inputs_payload_frame_line_pixel_2_0_11;
  assign inputsT_payload_frame_line_pixel_2_0_12 = inputs_payload_frame_line_pixel_2_0_12;
  assign inputsT_payload_frame_line_pixel_2_0_13 = inputs_payload_frame_line_pixel_2_0_13;
  assign inputsT_payload_frame_line_pixel_2_0_14 = inputs_payload_frame_line_pixel_2_0_14;
  assign inputsT_payload_frame_line_pixel_2_0_15 = inputs_payload_frame_line_pixel_2_0_15;
  assign inputsT_payload_frame_line_pixel_2_1_0 = inputs_payload_frame_line_pixel_2_1_0;
  assign inputsT_payload_frame_line_pixel_2_1_1 = inputs_payload_frame_line_pixel_2_1_1;
  assign inputsT_payload_frame_line_pixel_2_1_2 = inputs_payload_frame_line_pixel_2_1_2;
  assign inputsT_payload_frame_line_pixel_2_1_3 = inputs_payload_frame_line_pixel_2_1_3;
  assign inputsT_payload_frame_line_pixel_2_1_4 = inputs_payload_frame_line_pixel_2_1_4;
  assign inputsT_payload_frame_line_pixel_2_1_5 = inputs_payload_frame_line_pixel_2_1_5;
  assign inputsT_payload_frame_line_pixel_2_1_6 = inputs_payload_frame_line_pixel_2_1_6;
  assign inputsT_payload_frame_line_pixel_2_1_7 = inputs_payload_frame_line_pixel_2_1_7;
  assign inputsT_payload_frame_line_pixel_2_1_8 = inputs_payload_frame_line_pixel_2_1_8;
  assign inputsT_payload_frame_line_pixel_2_1_9 = inputs_payload_frame_line_pixel_2_1_9;
  assign inputsT_payload_frame_line_pixel_2_1_10 = inputs_payload_frame_line_pixel_2_1_10;
  assign inputsT_payload_frame_line_pixel_2_1_11 = inputs_payload_frame_line_pixel_2_1_11;
  assign inputsT_payload_frame_line_pixel_2_1_12 = inputs_payload_frame_line_pixel_2_1_12;
  assign inputsT_payload_frame_line_pixel_2_1_13 = inputs_payload_frame_line_pixel_2_1_13;
  assign inputsT_payload_frame_line_pixel_2_1_14 = inputs_payload_frame_line_pixel_2_1_14;
  assign inputsT_payload_frame_line_pixel_2_1_15 = inputs_payload_frame_line_pixel_2_1_15;
  assign inputsT_payload_frame_line_pixel_2_2_0 = inputs_payload_frame_line_pixel_2_2_0;
  assign inputsT_payload_frame_line_pixel_2_2_1 = inputs_payload_frame_line_pixel_2_2_1;
  assign inputsT_payload_frame_line_pixel_2_2_2 = inputs_payload_frame_line_pixel_2_2_2;
  assign inputsT_payload_frame_line_pixel_2_2_3 = inputs_payload_frame_line_pixel_2_2_3;
  assign inputsT_payload_frame_line_pixel_2_2_4 = inputs_payload_frame_line_pixel_2_2_4;
  assign inputsT_payload_frame_line_pixel_2_2_5 = inputs_payload_frame_line_pixel_2_2_5;
  assign inputsT_payload_frame_line_pixel_2_2_6 = inputs_payload_frame_line_pixel_2_2_6;
  assign inputsT_payload_frame_line_pixel_2_2_7 = inputs_payload_frame_line_pixel_2_2_7;
  assign inputsT_payload_frame_line_pixel_2_2_8 = inputs_payload_frame_line_pixel_2_2_8;
  assign inputsT_payload_frame_line_pixel_2_2_9 = inputs_payload_frame_line_pixel_2_2_9;
  assign inputsT_payload_frame_line_pixel_2_2_10 = inputs_payload_frame_line_pixel_2_2_10;
  assign inputsT_payload_frame_line_pixel_2_2_11 = inputs_payload_frame_line_pixel_2_2_11;
  assign inputsT_payload_frame_line_pixel_2_2_12 = inputs_payload_frame_line_pixel_2_2_12;
  assign inputsT_payload_frame_line_pixel_2_2_13 = inputs_payload_frame_line_pixel_2_2_13;
  assign inputsT_payload_frame_line_pixel_2_2_14 = inputs_payload_frame_line_pixel_2_2_14;
  assign inputsT_payload_frame_line_pixel_2_2_15 = inputs_payload_frame_line_pixel_2_2_15;
  assign inputsT_payload_frame_line_endOfLine = inputs_payload_frame_line_endOfLine;
  assign inputsT_payload_frame_endOfFrame = inputs_payload_frame_endOfFrame;
  assign inputsT_payload_endOfPack = inputs_payload_endOfPack;
  assign prevConv_valid = inputsT_valid;
  assign inputsT_ready = prevConv_ready;
  assign prevConv_payload_frame_line_pixel_0_0 = inputsT_payload_frame_line_pixel_0_0_0;
  assign prevConv_payload_frame_line_pixel_0_1 = weights_payload_0_0_0_0;
  assign prevConv_payload_frame_line_pixel_0_2 = weights_payload_1_0_0_0;
  assign prevConv_payload_frame_line_pixel_1_0 = inputsT_payload_frame_line_pixel_0_0_1;
  assign prevConv_payload_frame_line_pixel_1_1 = weights_payload_0_0_0_1;
  assign prevConv_payload_frame_line_pixel_1_2 = weights_payload_1_0_0_1;
  assign prevConv_payload_frame_line_pixel_2_0 = inputsT_payload_frame_line_pixel_0_0_2;
  assign prevConv_payload_frame_line_pixel_2_1 = weights_payload_0_0_0_2;
  assign prevConv_payload_frame_line_pixel_2_2 = weights_payload_1_0_0_2;
  assign prevConv_payload_frame_line_pixel_3_0 = inputsT_payload_frame_line_pixel_0_0_3;
  assign prevConv_payload_frame_line_pixel_3_1 = weights_payload_0_0_0_3;
  assign prevConv_payload_frame_line_pixel_3_2 = weights_payload_1_0_0_3;
  assign prevConv_payload_frame_line_pixel_4_0 = inputsT_payload_frame_line_pixel_0_0_4;
  assign prevConv_payload_frame_line_pixel_4_1 = weights_payload_0_0_0_4;
  assign prevConv_payload_frame_line_pixel_4_2 = weights_payload_1_0_0_4;
  assign prevConv_payload_frame_line_pixel_5_0 = inputsT_payload_frame_line_pixel_0_0_5;
  assign prevConv_payload_frame_line_pixel_5_1 = weights_payload_0_0_0_5;
  assign prevConv_payload_frame_line_pixel_5_2 = weights_payload_1_0_0_5;
  assign prevConv_payload_frame_line_pixel_6_0 = inputsT_payload_frame_line_pixel_0_0_6;
  assign prevConv_payload_frame_line_pixel_6_1 = weights_payload_0_0_0_6;
  assign prevConv_payload_frame_line_pixel_6_2 = weights_payload_1_0_0_6;
  assign prevConv_payload_frame_line_pixel_7_0 = inputsT_payload_frame_line_pixel_0_0_7;
  assign prevConv_payload_frame_line_pixel_7_1 = weights_payload_0_0_0_7;
  assign prevConv_payload_frame_line_pixel_7_2 = weights_payload_1_0_0_7;
  assign prevConv_payload_frame_line_pixel_8_0 = inputsT_payload_frame_line_pixel_0_0_8;
  assign prevConv_payload_frame_line_pixel_8_1 = weights_payload_0_0_0_8;
  assign prevConv_payload_frame_line_pixel_8_2 = weights_payload_1_0_0_8;
  assign prevConv_payload_frame_line_pixel_9_0 = inputsT_payload_frame_line_pixel_0_0_9;
  assign prevConv_payload_frame_line_pixel_9_1 = weights_payload_0_0_0_9;
  assign prevConv_payload_frame_line_pixel_9_2 = weights_payload_1_0_0_9;
  assign prevConv_payload_frame_line_pixel_10_0 = inputsT_payload_frame_line_pixel_0_0_10;
  assign prevConv_payload_frame_line_pixel_10_1 = weights_payload_0_0_0_10;
  assign prevConv_payload_frame_line_pixel_10_2 = weights_payload_1_0_0_10;
  assign prevConv_payload_frame_line_pixel_11_0 = inputsT_payload_frame_line_pixel_0_0_11;
  assign prevConv_payload_frame_line_pixel_11_1 = weights_payload_0_0_0_11;
  assign prevConv_payload_frame_line_pixel_11_2 = weights_payload_1_0_0_11;
  assign prevConv_payload_frame_line_pixel_12_0 = inputsT_payload_frame_line_pixel_0_0_12;
  assign prevConv_payload_frame_line_pixel_12_1 = weights_payload_0_0_0_12;
  assign prevConv_payload_frame_line_pixel_12_2 = weights_payload_1_0_0_12;
  assign prevConv_payload_frame_line_pixel_13_0 = inputsT_payload_frame_line_pixel_0_0_13;
  assign prevConv_payload_frame_line_pixel_13_1 = weights_payload_0_0_0_13;
  assign prevConv_payload_frame_line_pixel_13_2 = weights_payload_1_0_0_13;
  assign prevConv_payload_frame_line_pixel_14_0 = inputsT_payload_frame_line_pixel_0_0_14;
  assign prevConv_payload_frame_line_pixel_14_1 = weights_payload_0_0_0_14;
  assign prevConv_payload_frame_line_pixel_14_2 = weights_payload_1_0_0_14;
  assign prevConv_payload_frame_line_pixel_15_0 = inputsT_payload_frame_line_pixel_0_0_15;
  assign prevConv_payload_frame_line_pixel_15_1 = weights_payload_0_0_0_15;
  assign prevConv_payload_frame_line_pixel_15_2 = weights_payload_1_0_0_15;
  assign prevConv_payload_frame_line_pixel_16_0 = inputsT_payload_frame_line_pixel_0_1_0;
  assign prevConv_payload_frame_line_pixel_16_1 = weights_payload_0_0_1_0;
  assign prevConv_payload_frame_line_pixel_16_2 = weights_payload_1_0_1_0;
  assign prevConv_payload_frame_line_pixel_17_0 = inputsT_payload_frame_line_pixel_0_1_1;
  assign prevConv_payload_frame_line_pixel_17_1 = weights_payload_0_0_1_1;
  assign prevConv_payload_frame_line_pixel_17_2 = weights_payload_1_0_1_1;
  assign prevConv_payload_frame_line_pixel_18_0 = inputsT_payload_frame_line_pixel_0_1_2;
  assign prevConv_payload_frame_line_pixel_18_1 = weights_payload_0_0_1_2;
  assign prevConv_payload_frame_line_pixel_18_2 = weights_payload_1_0_1_2;
  assign prevConv_payload_frame_line_pixel_19_0 = inputsT_payload_frame_line_pixel_0_1_3;
  assign prevConv_payload_frame_line_pixel_19_1 = weights_payload_0_0_1_3;
  assign prevConv_payload_frame_line_pixel_19_2 = weights_payload_1_0_1_3;
  assign prevConv_payload_frame_line_pixel_20_0 = inputsT_payload_frame_line_pixel_0_1_4;
  assign prevConv_payload_frame_line_pixel_20_1 = weights_payload_0_0_1_4;
  assign prevConv_payload_frame_line_pixel_20_2 = weights_payload_1_0_1_4;
  assign prevConv_payload_frame_line_pixel_21_0 = inputsT_payload_frame_line_pixel_0_1_5;
  assign prevConv_payload_frame_line_pixel_21_1 = weights_payload_0_0_1_5;
  assign prevConv_payload_frame_line_pixel_21_2 = weights_payload_1_0_1_5;
  assign prevConv_payload_frame_line_pixel_22_0 = inputsT_payload_frame_line_pixel_0_1_6;
  assign prevConv_payload_frame_line_pixel_22_1 = weights_payload_0_0_1_6;
  assign prevConv_payload_frame_line_pixel_22_2 = weights_payload_1_0_1_6;
  assign prevConv_payload_frame_line_pixel_23_0 = inputsT_payload_frame_line_pixel_0_1_7;
  assign prevConv_payload_frame_line_pixel_23_1 = weights_payload_0_0_1_7;
  assign prevConv_payload_frame_line_pixel_23_2 = weights_payload_1_0_1_7;
  assign prevConv_payload_frame_line_pixel_24_0 = inputsT_payload_frame_line_pixel_0_1_8;
  assign prevConv_payload_frame_line_pixel_24_1 = weights_payload_0_0_1_8;
  assign prevConv_payload_frame_line_pixel_24_2 = weights_payload_1_0_1_8;
  assign prevConv_payload_frame_line_pixel_25_0 = inputsT_payload_frame_line_pixel_0_1_9;
  assign prevConv_payload_frame_line_pixel_25_1 = weights_payload_0_0_1_9;
  assign prevConv_payload_frame_line_pixel_25_2 = weights_payload_1_0_1_9;
  assign prevConv_payload_frame_line_pixel_26_0 = inputsT_payload_frame_line_pixel_0_1_10;
  assign prevConv_payload_frame_line_pixel_26_1 = weights_payload_0_0_1_10;
  assign prevConv_payload_frame_line_pixel_26_2 = weights_payload_1_0_1_10;
  assign prevConv_payload_frame_line_pixel_27_0 = inputsT_payload_frame_line_pixel_0_1_11;
  assign prevConv_payload_frame_line_pixel_27_1 = weights_payload_0_0_1_11;
  assign prevConv_payload_frame_line_pixel_27_2 = weights_payload_1_0_1_11;
  assign prevConv_payload_frame_line_pixel_28_0 = inputsT_payload_frame_line_pixel_0_1_12;
  assign prevConv_payload_frame_line_pixel_28_1 = weights_payload_0_0_1_12;
  assign prevConv_payload_frame_line_pixel_28_2 = weights_payload_1_0_1_12;
  assign prevConv_payload_frame_line_pixel_29_0 = inputsT_payload_frame_line_pixel_0_1_13;
  assign prevConv_payload_frame_line_pixel_29_1 = weights_payload_0_0_1_13;
  assign prevConv_payload_frame_line_pixel_29_2 = weights_payload_1_0_1_13;
  assign prevConv_payload_frame_line_pixel_30_0 = inputsT_payload_frame_line_pixel_0_1_14;
  assign prevConv_payload_frame_line_pixel_30_1 = weights_payload_0_0_1_14;
  assign prevConv_payload_frame_line_pixel_30_2 = weights_payload_1_0_1_14;
  assign prevConv_payload_frame_line_pixel_31_0 = inputsT_payload_frame_line_pixel_0_1_15;
  assign prevConv_payload_frame_line_pixel_31_1 = weights_payload_0_0_1_15;
  assign prevConv_payload_frame_line_pixel_31_2 = weights_payload_1_0_1_15;
  assign prevConv_payload_frame_line_pixel_32_0 = inputsT_payload_frame_line_pixel_0_2_0;
  assign prevConv_payload_frame_line_pixel_32_1 = weights_payload_0_0_2_0;
  assign prevConv_payload_frame_line_pixel_32_2 = weights_payload_1_0_2_0;
  assign prevConv_payload_frame_line_pixel_33_0 = inputsT_payload_frame_line_pixel_0_2_1;
  assign prevConv_payload_frame_line_pixel_33_1 = weights_payload_0_0_2_1;
  assign prevConv_payload_frame_line_pixel_33_2 = weights_payload_1_0_2_1;
  assign prevConv_payload_frame_line_pixel_34_0 = inputsT_payload_frame_line_pixel_0_2_2;
  assign prevConv_payload_frame_line_pixel_34_1 = weights_payload_0_0_2_2;
  assign prevConv_payload_frame_line_pixel_34_2 = weights_payload_1_0_2_2;
  assign prevConv_payload_frame_line_pixel_35_0 = inputsT_payload_frame_line_pixel_0_2_3;
  assign prevConv_payload_frame_line_pixel_35_1 = weights_payload_0_0_2_3;
  assign prevConv_payload_frame_line_pixel_35_2 = weights_payload_1_0_2_3;
  assign prevConv_payload_frame_line_pixel_36_0 = inputsT_payload_frame_line_pixel_0_2_4;
  assign prevConv_payload_frame_line_pixel_36_1 = weights_payload_0_0_2_4;
  assign prevConv_payload_frame_line_pixel_36_2 = weights_payload_1_0_2_4;
  assign prevConv_payload_frame_line_pixel_37_0 = inputsT_payload_frame_line_pixel_0_2_5;
  assign prevConv_payload_frame_line_pixel_37_1 = weights_payload_0_0_2_5;
  assign prevConv_payload_frame_line_pixel_37_2 = weights_payload_1_0_2_5;
  assign prevConv_payload_frame_line_pixel_38_0 = inputsT_payload_frame_line_pixel_0_2_6;
  assign prevConv_payload_frame_line_pixel_38_1 = weights_payload_0_0_2_6;
  assign prevConv_payload_frame_line_pixel_38_2 = weights_payload_1_0_2_6;
  assign prevConv_payload_frame_line_pixel_39_0 = inputsT_payload_frame_line_pixel_0_2_7;
  assign prevConv_payload_frame_line_pixel_39_1 = weights_payload_0_0_2_7;
  assign prevConv_payload_frame_line_pixel_39_2 = weights_payload_1_0_2_7;
  assign prevConv_payload_frame_line_pixel_40_0 = inputsT_payload_frame_line_pixel_0_2_8;
  assign prevConv_payload_frame_line_pixel_40_1 = weights_payload_0_0_2_8;
  assign prevConv_payload_frame_line_pixel_40_2 = weights_payload_1_0_2_8;
  assign prevConv_payload_frame_line_pixel_41_0 = inputsT_payload_frame_line_pixel_0_2_9;
  assign prevConv_payload_frame_line_pixel_41_1 = weights_payload_0_0_2_9;
  assign prevConv_payload_frame_line_pixel_41_2 = weights_payload_1_0_2_9;
  assign prevConv_payload_frame_line_pixel_42_0 = inputsT_payload_frame_line_pixel_0_2_10;
  assign prevConv_payload_frame_line_pixel_42_1 = weights_payload_0_0_2_10;
  assign prevConv_payload_frame_line_pixel_42_2 = weights_payload_1_0_2_10;
  assign prevConv_payload_frame_line_pixel_43_0 = inputsT_payload_frame_line_pixel_0_2_11;
  assign prevConv_payload_frame_line_pixel_43_1 = weights_payload_0_0_2_11;
  assign prevConv_payload_frame_line_pixel_43_2 = weights_payload_1_0_2_11;
  assign prevConv_payload_frame_line_pixel_44_0 = inputsT_payload_frame_line_pixel_0_2_12;
  assign prevConv_payload_frame_line_pixel_44_1 = weights_payload_0_0_2_12;
  assign prevConv_payload_frame_line_pixel_44_2 = weights_payload_1_0_2_12;
  assign prevConv_payload_frame_line_pixel_45_0 = inputsT_payload_frame_line_pixel_0_2_13;
  assign prevConv_payload_frame_line_pixel_45_1 = weights_payload_0_0_2_13;
  assign prevConv_payload_frame_line_pixel_45_2 = weights_payload_1_0_2_13;
  assign prevConv_payload_frame_line_pixel_46_0 = inputsT_payload_frame_line_pixel_0_2_14;
  assign prevConv_payload_frame_line_pixel_46_1 = weights_payload_0_0_2_14;
  assign prevConv_payload_frame_line_pixel_46_2 = weights_payload_1_0_2_14;
  assign prevConv_payload_frame_line_pixel_47_0 = inputsT_payload_frame_line_pixel_0_2_15;
  assign prevConv_payload_frame_line_pixel_47_1 = weights_payload_0_0_2_15;
  assign prevConv_payload_frame_line_pixel_47_2 = weights_payload_1_0_2_15;
  assign prevConv_payload_frame_line_pixel_48_0 = inputsT_payload_frame_line_pixel_1_0_0;
  assign prevConv_payload_frame_line_pixel_48_1 = weights_payload_0_1_0_0;
  assign prevConv_payload_frame_line_pixel_48_2 = weights_payload_1_1_0_0;
  assign prevConv_payload_frame_line_pixel_49_0 = inputsT_payload_frame_line_pixel_1_0_1;
  assign prevConv_payload_frame_line_pixel_49_1 = weights_payload_0_1_0_1;
  assign prevConv_payload_frame_line_pixel_49_2 = weights_payload_1_1_0_1;
  assign prevConv_payload_frame_line_pixel_50_0 = inputsT_payload_frame_line_pixel_1_0_2;
  assign prevConv_payload_frame_line_pixel_50_1 = weights_payload_0_1_0_2;
  assign prevConv_payload_frame_line_pixel_50_2 = weights_payload_1_1_0_2;
  assign prevConv_payload_frame_line_pixel_51_0 = inputsT_payload_frame_line_pixel_1_0_3;
  assign prevConv_payload_frame_line_pixel_51_1 = weights_payload_0_1_0_3;
  assign prevConv_payload_frame_line_pixel_51_2 = weights_payload_1_1_0_3;
  assign prevConv_payload_frame_line_pixel_52_0 = inputsT_payload_frame_line_pixel_1_0_4;
  assign prevConv_payload_frame_line_pixel_52_1 = weights_payload_0_1_0_4;
  assign prevConv_payload_frame_line_pixel_52_2 = weights_payload_1_1_0_4;
  assign prevConv_payload_frame_line_pixel_53_0 = inputsT_payload_frame_line_pixel_1_0_5;
  assign prevConv_payload_frame_line_pixel_53_1 = weights_payload_0_1_0_5;
  assign prevConv_payload_frame_line_pixel_53_2 = weights_payload_1_1_0_5;
  assign prevConv_payload_frame_line_pixel_54_0 = inputsT_payload_frame_line_pixel_1_0_6;
  assign prevConv_payload_frame_line_pixel_54_1 = weights_payload_0_1_0_6;
  assign prevConv_payload_frame_line_pixel_54_2 = weights_payload_1_1_0_6;
  assign prevConv_payload_frame_line_pixel_55_0 = inputsT_payload_frame_line_pixel_1_0_7;
  assign prevConv_payload_frame_line_pixel_55_1 = weights_payload_0_1_0_7;
  assign prevConv_payload_frame_line_pixel_55_2 = weights_payload_1_1_0_7;
  assign prevConv_payload_frame_line_pixel_56_0 = inputsT_payload_frame_line_pixel_1_0_8;
  assign prevConv_payload_frame_line_pixel_56_1 = weights_payload_0_1_0_8;
  assign prevConv_payload_frame_line_pixel_56_2 = weights_payload_1_1_0_8;
  assign prevConv_payload_frame_line_pixel_57_0 = inputsT_payload_frame_line_pixel_1_0_9;
  assign prevConv_payload_frame_line_pixel_57_1 = weights_payload_0_1_0_9;
  assign prevConv_payload_frame_line_pixel_57_2 = weights_payload_1_1_0_9;
  assign prevConv_payload_frame_line_pixel_58_0 = inputsT_payload_frame_line_pixel_1_0_10;
  assign prevConv_payload_frame_line_pixel_58_1 = weights_payload_0_1_0_10;
  assign prevConv_payload_frame_line_pixel_58_2 = weights_payload_1_1_0_10;
  assign prevConv_payload_frame_line_pixel_59_0 = inputsT_payload_frame_line_pixel_1_0_11;
  assign prevConv_payload_frame_line_pixel_59_1 = weights_payload_0_1_0_11;
  assign prevConv_payload_frame_line_pixel_59_2 = weights_payload_1_1_0_11;
  assign prevConv_payload_frame_line_pixel_60_0 = inputsT_payload_frame_line_pixel_1_0_12;
  assign prevConv_payload_frame_line_pixel_60_1 = weights_payload_0_1_0_12;
  assign prevConv_payload_frame_line_pixel_60_2 = weights_payload_1_1_0_12;
  assign prevConv_payload_frame_line_pixel_61_0 = inputsT_payload_frame_line_pixel_1_0_13;
  assign prevConv_payload_frame_line_pixel_61_1 = weights_payload_0_1_0_13;
  assign prevConv_payload_frame_line_pixel_61_2 = weights_payload_1_1_0_13;
  assign prevConv_payload_frame_line_pixel_62_0 = inputsT_payload_frame_line_pixel_1_0_14;
  assign prevConv_payload_frame_line_pixel_62_1 = weights_payload_0_1_0_14;
  assign prevConv_payload_frame_line_pixel_62_2 = weights_payload_1_1_0_14;
  assign prevConv_payload_frame_line_pixel_63_0 = inputsT_payload_frame_line_pixel_1_0_15;
  assign prevConv_payload_frame_line_pixel_63_1 = weights_payload_0_1_0_15;
  assign prevConv_payload_frame_line_pixel_63_2 = weights_payload_1_1_0_15;
  assign prevConv_payload_frame_line_pixel_64_0 = inputsT_payload_frame_line_pixel_1_1_0;
  assign prevConv_payload_frame_line_pixel_64_1 = weights_payload_0_1_1_0;
  assign prevConv_payload_frame_line_pixel_64_2 = weights_payload_1_1_1_0;
  assign prevConv_payload_frame_line_pixel_65_0 = inputsT_payload_frame_line_pixel_1_1_1;
  assign prevConv_payload_frame_line_pixel_65_1 = weights_payload_0_1_1_1;
  assign prevConv_payload_frame_line_pixel_65_2 = weights_payload_1_1_1_1;
  assign prevConv_payload_frame_line_pixel_66_0 = inputsT_payload_frame_line_pixel_1_1_2;
  assign prevConv_payload_frame_line_pixel_66_1 = weights_payload_0_1_1_2;
  assign prevConv_payload_frame_line_pixel_66_2 = weights_payload_1_1_1_2;
  assign prevConv_payload_frame_line_pixel_67_0 = inputsT_payload_frame_line_pixel_1_1_3;
  assign prevConv_payload_frame_line_pixel_67_1 = weights_payload_0_1_1_3;
  assign prevConv_payload_frame_line_pixel_67_2 = weights_payload_1_1_1_3;
  assign prevConv_payload_frame_line_pixel_68_0 = inputsT_payload_frame_line_pixel_1_1_4;
  assign prevConv_payload_frame_line_pixel_68_1 = weights_payload_0_1_1_4;
  assign prevConv_payload_frame_line_pixel_68_2 = weights_payload_1_1_1_4;
  assign prevConv_payload_frame_line_pixel_69_0 = inputsT_payload_frame_line_pixel_1_1_5;
  assign prevConv_payload_frame_line_pixel_69_1 = weights_payload_0_1_1_5;
  assign prevConv_payload_frame_line_pixel_69_2 = weights_payload_1_1_1_5;
  assign prevConv_payload_frame_line_pixel_70_0 = inputsT_payload_frame_line_pixel_1_1_6;
  assign prevConv_payload_frame_line_pixel_70_1 = weights_payload_0_1_1_6;
  assign prevConv_payload_frame_line_pixel_70_2 = weights_payload_1_1_1_6;
  assign prevConv_payload_frame_line_pixel_71_0 = inputsT_payload_frame_line_pixel_1_1_7;
  assign prevConv_payload_frame_line_pixel_71_1 = weights_payload_0_1_1_7;
  assign prevConv_payload_frame_line_pixel_71_2 = weights_payload_1_1_1_7;
  assign prevConv_payload_frame_line_pixel_72_0 = inputsT_payload_frame_line_pixel_1_1_8;
  assign prevConv_payload_frame_line_pixel_72_1 = weights_payload_0_1_1_8;
  assign prevConv_payload_frame_line_pixel_72_2 = weights_payload_1_1_1_8;
  assign prevConv_payload_frame_line_pixel_73_0 = inputsT_payload_frame_line_pixel_1_1_9;
  assign prevConv_payload_frame_line_pixel_73_1 = weights_payload_0_1_1_9;
  assign prevConv_payload_frame_line_pixel_73_2 = weights_payload_1_1_1_9;
  assign prevConv_payload_frame_line_pixel_74_0 = inputsT_payload_frame_line_pixel_1_1_10;
  assign prevConv_payload_frame_line_pixel_74_1 = weights_payload_0_1_1_10;
  assign prevConv_payload_frame_line_pixel_74_2 = weights_payload_1_1_1_10;
  assign prevConv_payload_frame_line_pixel_75_0 = inputsT_payload_frame_line_pixel_1_1_11;
  assign prevConv_payload_frame_line_pixel_75_1 = weights_payload_0_1_1_11;
  assign prevConv_payload_frame_line_pixel_75_2 = weights_payload_1_1_1_11;
  assign prevConv_payload_frame_line_pixel_76_0 = inputsT_payload_frame_line_pixel_1_1_12;
  assign prevConv_payload_frame_line_pixel_76_1 = weights_payload_0_1_1_12;
  assign prevConv_payload_frame_line_pixel_76_2 = weights_payload_1_1_1_12;
  assign prevConv_payload_frame_line_pixel_77_0 = inputsT_payload_frame_line_pixel_1_1_13;
  assign prevConv_payload_frame_line_pixel_77_1 = weights_payload_0_1_1_13;
  assign prevConv_payload_frame_line_pixel_77_2 = weights_payload_1_1_1_13;
  assign prevConv_payload_frame_line_pixel_78_0 = inputsT_payload_frame_line_pixel_1_1_14;
  assign prevConv_payload_frame_line_pixel_78_1 = weights_payload_0_1_1_14;
  assign prevConv_payload_frame_line_pixel_78_2 = weights_payload_1_1_1_14;
  assign prevConv_payload_frame_line_pixel_79_0 = inputsT_payload_frame_line_pixel_1_1_15;
  assign prevConv_payload_frame_line_pixel_79_1 = weights_payload_0_1_1_15;
  assign prevConv_payload_frame_line_pixel_79_2 = weights_payload_1_1_1_15;
  assign prevConv_payload_frame_line_pixel_80_0 = inputsT_payload_frame_line_pixel_1_2_0;
  assign prevConv_payload_frame_line_pixel_80_1 = weights_payload_0_1_2_0;
  assign prevConv_payload_frame_line_pixel_80_2 = weights_payload_1_1_2_0;
  assign prevConv_payload_frame_line_pixel_81_0 = inputsT_payload_frame_line_pixel_1_2_1;
  assign prevConv_payload_frame_line_pixel_81_1 = weights_payload_0_1_2_1;
  assign prevConv_payload_frame_line_pixel_81_2 = weights_payload_1_1_2_1;
  assign prevConv_payload_frame_line_pixel_82_0 = inputsT_payload_frame_line_pixel_1_2_2;
  assign prevConv_payload_frame_line_pixel_82_1 = weights_payload_0_1_2_2;
  assign prevConv_payload_frame_line_pixel_82_2 = weights_payload_1_1_2_2;
  assign prevConv_payload_frame_line_pixel_83_0 = inputsT_payload_frame_line_pixel_1_2_3;
  assign prevConv_payload_frame_line_pixel_83_1 = weights_payload_0_1_2_3;
  assign prevConv_payload_frame_line_pixel_83_2 = weights_payload_1_1_2_3;
  assign prevConv_payload_frame_line_pixel_84_0 = inputsT_payload_frame_line_pixel_1_2_4;
  assign prevConv_payload_frame_line_pixel_84_1 = weights_payload_0_1_2_4;
  assign prevConv_payload_frame_line_pixel_84_2 = weights_payload_1_1_2_4;
  assign prevConv_payload_frame_line_pixel_85_0 = inputsT_payload_frame_line_pixel_1_2_5;
  assign prevConv_payload_frame_line_pixel_85_1 = weights_payload_0_1_2_5;
  assign prevConv_payload_frame_line_pixel_85_2 = weights_payload_1_1_2_5;
  assign prevConv_payload_frame_line_pixel_86_0 = inputsT_payload_frame_line_pixel_1_2_6;
  assign prevConv_payload_frame_line_pixel_86_1 = weights_payload_0_1_2_6;
  assign prevConv_payload_frame_line_pixel_86_2 = weights_payload_1_1_2_6;
  assign prevConv_payload_frame_line_pixel_87_0 = inputsT_payload_frame_line_pixel_1_2_7;
  assign prevConv_payload_frame_line_pixel_87_1 = weights_payload_0_1_2_7;
  assign prevConv_payload_frame_line_pixel_87_2 = weights_payload_1_1_2_7;
  assign prevConv_payload_frame_line_pixel_88_0 = inputsT_payload_frame_line_pixel_1_2_8;
  assign prevConv_payload_frame_line_pixel_88_1 = weights_payload_0_1_2_8;
  assign prevConv_payload_frame_line_pixel_88_2 = weights_payload_1_1_2_8;
  assign prevConv_payload_frame_line_pixel_89_0 = inputsT_payload_frame_line_pixel_1_2_9;
  assign prevConv_payload_frame_line_pixel_89_1 = weights_payload_0_1_2_9;
  assign prevConv_payload_frame_line_pixel_89_2 = weights_payload_1_1_2_9;
  assign prevConv_payload_frame_line_pixel_90_0 = inputsT_payload_frame_line_pixel_1_2_10;
  assign prevConv_payload_frame_line_pixel_90_1 = weights_payload_0_1_2_10;
  assign prevConv_payload_frame_line_pixel_90_2 = weights_payload_1_1_2_10;
  assign prevConv_payload_frame_line_pixel_91_0 = inputsT_payload_frame_line_pixel_1_2_11;
  assign prevConv_payload_frame_line_pixel_91_1 = weights_payload_0_1_2_11;
  assign prevConv_payload_frame_line_pixel_91_2 = weights_payload_1_1_2_11;
  assign prevConv_payload_frame_line_pixel_92_0 = inputsT_payload_frame_line_pixel_1_2_12;
  assign prevConv_payload_frame_line_pixel_92_1 = weights_payload_0_1_2_12;
  assign prevConv_payload_frame_line_pixel_92_2 = weights_payload_1_1_2_12;
  assign prevConv_payload_frame_line_pixel_93_0 = inputsT_payload_frame_line_pixel_1_2_13;
  assign prevConv_payload_frame_line_pixel_93_1 = weights_payload_0_1_2_13;
  assign prevConv_payload_frame_line_pixel_93_2 = weights_payload_1_1_2_13;
  assign prevConv_payload_frame_line_pixel_94_0 = inputsT_payload_frame_line_pixel_1_2_14;
  assign prevConv_payload_frame_line_pixel_94_1 = weights_payload_0_1_2_14;
  assign prevConv_payload_frame_line_pixel_94_2 = weights_payload_1_1_2_14;
  assign prevConv_payload_frame_line_pixel_95_0 = inputsT_payload_frame_line_pixel_1_2_15;
  assign prevConv_payload_frame_line_pixel_95_1 = weights_payload_0_1_2_15;
  assign prevConv_payload_frame_line_pixel_95_2 = weights_payload_1_1_2_15;
  assign prevConv_payload_frame_line_pixel_96_0 = inputsT_payload_frame_line_pixel_2_0_0;
  assign prevConv_payload_frame_line_pixel_96_1 = weights_payload_0_2_0_0;
  assign prevConv_payload_frame_line_pixel_96_2 = weights_payload_1_2_0_0;
  assign prevConv_payload_frame_line_pixel_97_0 = inputsT_payload_frame_line_pixel_2_0_1;
  assign prevConv_payload_frame_line_pixel_97_1 = weights_payload_0_2_0_1;
  assign prevConv_payload_frame_line_pixel_97_2 = weights_payload_1_2_0_1;
  assign prevConv_payload_frame_line_pixel_98_0 = inputsT_payload_frame_line_pixel_2_0_2;
  assign prevConv_payload_frame_line_pixel_98_1 = weights_payload_0_2_0_2;
  assign prevConv_payload_frame_line_pixel_98_2 = weights_payload_1_2_0_2;
  assign prevConv_payload_frame_line_pixel_99_0 = inputsT_payload_frame_line_pixel_2_0_3;
  assign prevConv_payload_frame_line_pixel_99_1 = weights_payload_0_2_0_3;
  assign prevConv_payload_frame_line_pixel_99_2 = weights_payload_1_2_0_3;
  assign prevConv_payload_frame_line_pixel_100_0 = inputsT_payload_frame_line_pixel_2_0_4;
  assign prevConv_payload_frame_line_pixel_100_1 = weights_payload_0_2_0_4;
  assign prevConv_payload_frame_line_pixel_100_2 = weights_payload_1_2_0_4;
  assign prevConv_payload_frame_line_pixel_101_0 = inputsT_payload_frame_line_pixel_2_0_5;
  assign prevConv_payload_frame_line_pixel_101_1 = weights_payload_0_2_0_5;
  assign prevConv_payload_frame_line_pixel_101_2 = weights_payload_1_2_0_5;
  assign prevConv_payload_frame_line_pixel_102_0 = inputsT_payload_frame_line_pixel_2_0_6;
  assign prevConv_payload_frame_line_pixel_102_1 = weights_payload_0_2_0_6;
  assign prevConv_payload_frame_line_pixel_102_2 = weights_payload_1_2_0_6;
  assign prevConv_payload_frame_line_pixel_103_0 = inputsT_payload_frame_line_pixel_2_0_7;
  assign prevConv_payload_frame_line_pixel_103_1 = weights_payload_0_2_0_7;
  assign prevConv_payload_frame_line_pixel_103_2 = weights_payload_1_2_0_7;
  assign prevConv_payload_frame_line_pixel_104_0 = inputsT_payload_frame_line_pixel_2_0_8;
  assign prevConv_payload_frame_line_pixel_104_1 = weights_payload_0_2_0_8;
  assign prevConv_payload_frame_line_pixel_104_2 = weights_payload_1_2_0_8;
  assign prevConv_payload_frame_line_pixel_105_0 = inputsT_payload_frame_line_pixel_2_0_9;
  assign prevConv_payload_frame_line_pixel_105_1 = weights_payload_0_2_0_9;
  assign prevConv_payload_frame_line_pixel_105_2 = weights_payload_1_2_0_9;
  assign prevConv_payload_frame_line_pixel_106_0 = inputsT_payload_frame_line_pixel_2_0_10;
  assign prevConv_payload_frame_line_pixel_106_1 = weights_payload_0_2_0_10;
  assign prevConv_payload_frame_line_pixel_106_2 = weights_payload_1_2_0_10;
  assign prevConv_payload_frame_line_pixel_107_0 = inputsT_payload_frame_line_pixel_2_0_11;
  assign prevConv_payload_frame_line_pixel_107_1 = weights_payload_0_2_0_11;
  assign prevConv_payload_frame_line_pixel_107_2 = weights_payload_1_2_0_11;
  assign prevConv_payload_frame_line_pixel_108_0 = inputsT_payload_frame_line_pixel_2_0_12;
  assign prevConv_payload_frame_line_pixel_108_1 = weights_payload_0_2_0_12;
  assign prevConv_payload_frame_line_pixel_108_2 = weights_payload_1_2_0_12;
  assign prevConv_payload_frame_line_pixel_109_0 = inputsT_payload_frame_line_pixel_2_0_13;
  assign prevConv_payload_frame_line_pixel_109_1 = weights_payload_0_2_0_13;
  assign prevConv_payload_frame_line_pixel_109_2 = weights_payload_1_2_0_13;
  assign prevConv_payload_frame_line_pixel_110_0 = inputsT_payload_frame_line_pixel_2_0_14;
  assign prevConv_payload_frame_line_pixel_110_1 = weights_payload_0_2_0_14;
  assign prevConv_payload_frame_line_pixel_110_2 = weights_payload_1_2_0_14;
  assign prevConv_payload_frame_line_pixel_111_0 = inputsT_payload_frame_line_pixel_2_0_15;
  assign prevConv_payload_frame_line_pixel_111_1 = weights_payload_0_2_0_15;
  assign prevConv_payload_frame_line_pixel_111_2 = weights_payload_1_2_0_15;
  assign prevConv_payload_frame_line_pixel_112_0 = inputsT_payload_frame_line_pixel_2_1_0;
  assign prevConv_payload_frame_line_pixel_112_1 = weights_payload_0_2_1_0;
  assign prevConv_payload_frame_line_pixel_112_2 = weights_payload_1_2_1_0;
  assign prevConv_payload_frame_line_pixel_113_0 = inputsT_payload_frame_line_pixel_2_1_1;
  assign prevConv_payload_frame_line_pixel_113_1 = weights_payload_0_2_1_1;
  assign prevConv_payload_frame_line_pixel_113_2 = weights_payload_1_2_1_1;
  assign prevConv_payload_frame_line_pixel_114_0 = inputsT_payload_frame_line_pixel_2_1_2;
  assign prevConv_payload_frame_line_pixel_114_1 = weights_payload_0_2_1_2;
  assign prevConv_payload_frame_line_pixel_114_2 = weights_payload_1_2_1_2;
  assign prevConv_payload_frame_line_pixel_115_0 = inputsT_payload_frame_line_pixel_2_1_3;
  assign prevConv_payload_frame_line_pixel_115_1 = weights_payload_0_2_1_3;
  assign prevConv_payload_frame_line_pixel_115_2 = weights_payload_1_2_1_3;
  assign prevConv_payload_frame_line_pixel_116_0 = inputsT_payload_frame_line_pixel_2_1_4;
  assign prevConv_payload_frame_line_pixel_116_1 = weights_payload_0_2_1_4;
  assign prevConv_payload_frame_line_pixel_116_2 = weights_payload_1_2_1_4;
  assign prevConv_payload_frame_line_pixel_117_0 = inputsT_payload_frame_line_pixel_2_1_5;
  assign prevConv_payload_frame_line_pixel_117_1 = weights_payload_0_2_1_5;
  assign prevConv_payload_frame_line_pixel_117_2 = weights_payload_1_2_1_5;
  assign prevConv_payload_frame_line_pixel_118_0 = inputsT_payload_frame_line_pixel_2_1_6;
  assign prevConv_payload_frame_line_pixel_118_1 = weights_payload_0_2_1_6;
  assign prevConv_payload_frame_line_pixel_118_2 = weights_payload_1_2_1_6;
  assign prevConv_payload_frame_line_pixel_119_0 = inputsT_payload_frame_line_pixel_2_1_7;
  assign prevConv_payload_frame_line_pixel_119_1 = weights_payload_0_2_1_7;
  assign prevConv_payload_frame_line_pixel_119_2 = weights_payload_1_2_1_7;
  assign prevConv_payload_frame_line_pixel_120_0 = inputsT_payload_frame_line_pixel_2_1_8;
  assign prevConv_payload_frame_line_pixel_120_1 = weights_payload_0_2_1_8;
  assign prevConv_payload_frame_line_pixel_120_2 = weights_payload_1_2_1_8;
  assign prevConv_payload_frame_line_pixel_121_0 = inputsT_payload_frame_line_pixel_2_1_9;
  assign prevConv_payload_frame_line_pixel_121_1 = weights_payload_0_2_1_9;
  assign prevConv_payload_frame_line_pixel_121_2 = weights_payload_1_2_1_9;
  assign prevConv_payload_frame_line_pixel_122_0 = inputsT_payload_frame_line_pixel_2_1_10;
  assign prevConv_payload_frame_line_pixel_122_1 = weights_payload_0_2_1_10;
  assign prevConv_payload_frame_line_pixel_122_2 = weights_payload_1_2_1_10;
  assign prevConv_payload_frame_line_pixel_123_0 = inputsT_payload_frame_line_pixel_2_1_11;
  assign prevConv_payload_frame_line_pixel_123_1 = weights_payload_0_2_1_11;
  assign prevConv_payload_frame_line_pixel_123_2 = weights_payload_1_2_1_11;
  assign prevConv_payload_frame_line_pixel_124_0 = inputsT_payload_frame_line_pixel_2_1_12;
  assign prevConv_payload_frame_line_pixel_124_1 = weights_payload_0_2_1_12;
  assign prevConv_payload_frame_line_pixel_124_2 = weights_payload_1_2_1_12;
  assign prevConv_payload_frame_line_pixel_125_0 = inputsT_payload_frame_line_pixel_2_1_13;
  assign prevConv_payload_frame_line_pixel_125_1 = weights_payload_0_2_1_13;
  assign prevConv_payload_frame_line_pixel_125_2 = weights_payload_1_2_1_13;
  assign prevConv_payload_frame_line_pixel_126_0 = inputsT_payload_frame_line_pixel_2_1_14;
  assign prevConv_payload_frame_line_pixel_126_1 = weights_payload_0_2_1_14;
  assign prevConv_payload_frame_line_pixel_126_2 = weights_payload_1_2_1_14;
  assign prevConv_payload_frame_line_pixel_127_0 = inputsT_payload_frame_line_pixel_2_1_15;
  assign prevConv_payload_frame_line_pixel_127_1 = weights_payload_0_2_1_15;
  assign prevConv_payload_frame_line_pixel_127_2 = weights_payload_1_2_1_15;
  assign prevConv_payload_frame_line_pixel_128_0 = inputsT_payload_frame_line_pixel_2_2_0;
  assign prevConv_payload_frame_line_pixel_128_1 = weights_payload_0_2_2_0;
  assign prevConv_payload_frame_line_pixel_128_2 = weights_payload_1_2_2_0;
  assign prevConv_payload_frame_line_pixel_129_0 = inputsT_payload_frame_line_pixel_2_2_1;
  assign prevConv_payload_frame_line_pixel_129_1 = weights_payload_0_2_2_1;
  assign prevConv_payload_frame_line_pixel_129_2 = weights_payload_1_2_2_1;
  assign prevConv_payload_frame_line_pixel_130_0 = inputsT_payload_frame_line_pixel_2_2_2;
  assign prevConv_payload_frame_line_pixel_130_1 = weights_payload_0_2_2_2;
  assign prevConv_payload_frame_line_pixel_130_2 = weights_payload_1_2_2_2;
  assign prevConv_payload_frame_line_pixel_131_0 = inputsT_payload_frame_line_pixel_2_2_3;
  assign prevConv_payload_frame_line_pixel_131_1 = weights_payload_0_2_2_3;
  assign prevConv_payload_frame_line_pixel_131_2 = weights_payload_1_2_2_3;
  assign prevConv_payload_frame_line_pixel_132_0 = inputsT_payload_frame_line_pixel_2_2_4;
  assign prevConv_payload_frame_line_pixel_132_1 = weights_payload_0_2_2_4;
  assign prevConv_payload_frame_line_pixel_132_2 = weights_payload_1_2_2_4;
  assign prevConv_payload_frame_line_pixel_133_0 = inputsT_payload_frame_line_pixel_2_2_5;
  assign prevConv_payload_frame_line_pixel_133_1 = weights_payload_0_2_2_5;
  assign prevConv_payload_frame_line_pixel_133_2 = weights_payload_1_2_2_5;
  assign prevConv_payload_frame_line_pixel_134_0 = inputsT_payload_frame_line_pixel_2_2_6;
  assign prevConv_payload_frame_line_pixel_134_1 = weights_payload_0_2_2_6;
  assign prevConv_payload_frame_line_pixel_134_2 = weights_payload_1_2_2_6;
  assign prevConv_payload_frame_line_pixel_135_0 = inputsT_payload_frame_line_pixel_2_2_7;
  assign prevConv_payload_frame_line_pixel_135_1 = weights_payload_0_2_2_7;
  assign prevConv_payload_frame_line_pixel_135_2 = weights_payload_1_2_2_7;
  assign prevConv_payload_frame_line_pixel_136_0 = inputsT_payload_frame_line_pixel_2_2_8;
  assign prevConv_payload_frame_line_pixel_136_1 = weights_payload_0_2_2_8;
  assign prevConv_payload_frame_line_pixel_136_2 = weights_payload_1_2_2_8;
  assign prevConv_payload_frame_line_pixel_137_0 = inputsT_payload_frame_line_pixel_2_2_9;
  assign prevConv_payload_frame_line_pixel_137_1 = weights_payload_0_2_2_9;
  assign prevConv_payload_frame_line_pixel_137_2 = weights_payload_1_2_2_9;
  assign prevConv_payload_frame_line_pixel_138_0 = inputsT_payload_frame_line_pixel_2_2_10;
  assign prevConv_payload_frame_line_pixel_138_1 = weights_payload_0_2_2_10;
  assign prevConv_payload_frame_line_pixel_138_2 = weights_payload_1_2_2_10;
  assign prevConv_payload_frame_line_pixel_139_0 = inputsT_payload_frame_line_pixel_2_2_11;
  assign prevConv_payload_frame_line_pixel_139_1 = weights_payload_0_2_2_11;
  assign prevConv_payload_frame_line_pixel_139_2 = weights_payload_1_2_2_11;
  assign prevConv_payload_frame_line_pixel_140_0 = inputsT_payload_frame_line_pixel_2_2_12;
  assign prevConv_payload_frame_line_pixel_140_1 = weights_payload_0_2_2_12;
  assign prevConv_payload_frame_line_pixel_140_2 = weights_payload_1_2_2_12;
  assign prevConv_payload_frame_line_pixel_141_0 = inputsT_payload_frame_line_pixel_2_2_13;
  assign prevConv_payload_frame_line_pixel_141_1 = weights_payload_0_2_2_13;
  assign prevConv_payload_frame_line_pixel_141_2 = weights_payload_1_2_2_13;
  assign prevConv_payload_frame_line_pixel_142_0 = inputsT_payload_frame_line_pixel_2_2_14;
  assign prevConv_payload_frame_line_pixel_142_1 = weights_payload_0_2_2_14;
  assign prevConv_payload_frame_line_pixel_142_2 = weights_payload_1_2_2_14;
  assign prevConv_payload_frame_line_pixel_143_0 = inputsT_payload_frame_line_pixel_2_2_15;
  assign prevConv_payload_frame_line_pixel_143_1 = weights_payload_0_2_2_15;
  assign prevConv_payload_frame_line_pixel_143_2 = weights_payload_1_2_2_15;
  assign prevConv_payload_frame_line_endOfLine = inputsT_payload_frame_line_endOfLine;
  assign prevConv_payload_frame_endOfFrame = inputsT_payload_frame_endOfFrame;
  assign prevConv_payload_endOfPack = inputsT_payload_endOfPack;
  assign prevConv_ready = eventM2sPipes_9_eventIn_ready;
  assign postConv_payload_frame_line_pixel_0 = tmp_postConv_payload_frame_line_pixel_0_72;
  assign postConv_payload_frame_line_pixel_1 = tmp_postConv_payload_frame_line_pixel_1_72;
  assign postConv_valid = eventM2sPipes_9_eventOut_valid;
  assign postConv_payload_endOfPack = tmp_postConv_payload_endOfPack_8;
  assign postConv_payload_frame_endOfFrame = tmp_postConv_payload_frame_endOfFrame_8;
  assign postConv_payload_frame_line_endOfLine = tmp_postConv_payload_frame_line_endOfLine_8;
  assign inputsT_fire = (inputsT_valid && inputsT_ready);
  assign weights_ready = (inputsT_fire && inputsT_payload_frame_endOfFrame);
  assign postConv_ready = (! postConv_rValid);
  assign postConv_s2mPipe_valid = (postConv_valid || postConv_rValid);
  assign postConv_s2mPipe_payload_frame_line_pixel_0 = (postConv_rValid ? postConv_rData_frame_line_pixel_0 : postConv_payload_frame_line_pixel_0);
  assign postConv_s2mPipe_payload_frame_line_pixel_1 = (postConv_rValid ? postConv_rData_frame_line_pixel_1 : postConv_payload_frame_line_pixel_1);
  assign postConv_s2mPipe_payload_frame_line_endOfLine = (postConv_rValid ? postConv_rData_frame_line_endOfLine : postConv_payload_frame_line_endOfLine);
  assign postConv_s2mPipe_payload_frame_endOfFrame = (postConv_rValid ? postConv_rData_frame_endOfFrame : postConv_payload_frame_endOfFrame);
  assign postConv_s2mPipe_payload_endOfPack = (postConv_rValid ? postConv_rData_endOfPack : postConv_payload_endOfPack);
  assign postConv_s2mPipe_ready = acc_videoIn_ready;
  assign outputs_valid = acc_videoOut_valid;
  assign outputs_payload_frame_line_pixel_0 = acc_videoOut_payload_frame_line_pixel_0;
  assign outputs_payload_frame_line_pixel_1 = acc_videoOut_payload_frame_line_pixel_1;
  assign outputs_payload_frame_line_endOfLine = acc_videoOut_payload_frame_line_endOfLine;
  assign outputs_payload_frame_endOfFrame = acc_videoOut_payload_frame_endOfFrame;
  assign outputs_payload_endOfPack = acc_videoOut_payload_endOfPack;
  always @(posedge clk) begin
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0) + $signed(sIMD2INT8_1154_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_1 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_1) + $signed(sIMD2INT8_1157_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_2 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_2) + $signed(sIMD2INT8_1160_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_3 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_3) + $signed(sIMD2INT8_1163_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_4 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_4) + $signed(sIMD2INT8_1166_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_5 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_5) + $signed(sIMD2INT8_1169_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_6 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_6) + $signed(sIMD2INT8_1172_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_7 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_7) + $signed(sIMD2INT8_1175_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_8 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_8) + $signed(sIMD2INT8_1178_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_9 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_9) + $signed(sIMD2INT8_1181_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_10 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_10) + $signed(sIMD2INT8_1184_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_11 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_11) + $signed(sIMD2INT8_1187_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_12 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_12) + $signed(sIMD2INT8_1190_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_13 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_13) + $signed(sIMD2INT8_1193_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_14 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_14) + $signed(sIMD2INT8_1196_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_15 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_15) + $signed(sIMD2INT8_1199_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_16 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_16) + $signed(sIMD2INT8_1202_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_17 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_17) + $signed(sIMD2INT8_1205_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_18 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_18) + $signed(sIMD2INT8_1208_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_19 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_19) + $signed(sIMD2INT8_1211_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_20 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_20) + $signed(sIMD2INT8_1214_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_21 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_21) + $signed(sIMD2INT8_1217_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_22 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_22) + $signed(sIMD2INT8_1220_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_23 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_23) + $signed(sIMD2INT8_1223_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_24 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_24) + $signed(sIMD2INT8_1226_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_25 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_25) + $signed(sIMD2INT8_1229_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_26 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_26) + $signed(sIMD2INT8_1232_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_27 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_27) + $signed(sIMD2INT8_1235_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_28 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_28) + $signed(sIMD2INT8_1238_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_29 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_29) + $signed(sIMD2INT8_1241_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_30 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_30) + $signed(sIMD2INT8_1244_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_31 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_31) + $signed(sIMD2INT8_1247_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_32 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_32) + $signed(sIMD2INT8_1250_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_33 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_33) + $signed(sIMD2INT8_1253_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_34 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_34) + $signed(sIMD2INT8_1256_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_35 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_35) + $signed(sIMD2INT8_1259_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_36 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_36) + $signed(sIMD2INT8_1262_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_37 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_37) + $signed(sIMD2INT8_1265_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_38 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_38) + $signed(sIMD2INT8_1268_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_39 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_39) + $signed(sIMD2INT8_1271_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_40 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_40) + $signed(sIMD2INT8_1274_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_41 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_41) + $signed(sIMD2INT8_1277_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_42 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_42) + $signed(sIMD2INT8_1280_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_43 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_43) + $signed(sIMD2INT8_1283_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_44 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_44) + $signed(sIMD2INT8_1286_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_45 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_45) + $signed(sIMD2INT8_1289_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_46 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_46) + $signed(sIMD2INT8_1292_ab));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_0_47 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_47) + $signed(sIMD2INT8_1295_ab));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_48 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_48) + $signed(tmp_postConv_payload_frame_line_pixel_0_2));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_49 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_49) + $signed(tmp_postConv_payload_frame_line_pixel_0_5));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_50 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_50) + $signed(tmp_postConv_payload_frame_line_pixel_0_8));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_51 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_51) + $signed(tmp_postConv_payload_frame_line_pixel_0_11));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_52 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_52) + $signed(tmp_postConv_payload_frame_line_pixel_0_14));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_53 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_53) + $signed(tmp_postConv_payload_frame_line_pixel_0_17));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_54 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_54) + $signed(tmp_postConv_payload_frame_line_pixel_0_20));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_55 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_55) + $signed(tmp_postConv_payload_frame_line_pixel_0_23));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_56 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_56) + $signed(tmp_postConv_payload_frame_line_pixel_0_26));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_57 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_57) + $signed(tmp_postConv_payload_frame_line_pixel_0_29));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_58 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_58) + $signed(tmp_postConv_payload_frame_line_pixel_0_32));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_59 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_59) + $signed(tmp_postConv_payload_frame_line_pixel_0_35));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_60 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_60) + $signed(tmp_postConv_payload_frame_line_pixel_0_38));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_61 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_61) + $signed(tmp_postConv_payload_frame_line_pixel_0_41));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_62 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_62) + $signed(tmp_postConv_payload_frame_line_pixel_0_44));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_0_63 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_63) + $signed(tmp_postConv_payload_frame_line_pixel_0_47));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_64 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_64) + $signed(tmp_postConv_payload_frame_line_pixel_0_50));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_65 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_65) + $signed(tmp_postConv_payload_frame_line_pixel_0_53));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_66 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_66) + $signed(tmp_postConv_payload_frame_line_pixel_0_56));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_67 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_67) + $signed(tmp_postConv_payload_frame_line_pixel_0_59));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_68 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_68) + $signed(tmp_postConv_payload_frame_line_pixel_0_62));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_0_69 <= tmp_postConv_payload_frame_line_pixel_0_63;
    end
    if(eventM2sPipes_9_CEs_7) begin
      tmp_postConv_payload_frame_line_pixel_0_70 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_70) + $signed(tmp_postConv_payload_frame_line_pixel_0_66));
    end
    if(eventM2sPipes_9_CEs_7) begin
      tmp_postConv_payload_frame_line_pixel_0_71 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_71) + $signed(tmp_postConv_payload_frame_line_pixel_0_69));
    end
    if(eventM2sPipes_9_CEs_8) begin
      tmp_postConv_payload_frame_line_pixel_0_72 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_0_72) + $signed(tmp_tmp_postConv_payload_frame_line_pixel_0_72_1));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1) + $signed(sIMD2INT8_1154_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_1 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_1) + $signed(sIMD2INT8_1157_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_2 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_2) + $signed(sIMD2INT8_1160_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_3 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_3) + $signed(sIMD2INT8_1163_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_4 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_4) + $signed(sIMD2INT8_1166_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_5 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_5) + $signed(sIMD2INT8_1169_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_6 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_6) + $signed(sIMD2INT8_1172_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_7 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_7) + $signed(sIMD2INT8_1175_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_8 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_8) + $signed(sIMD2INT8_1178_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_9 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_9) + $signed(sIMD2INT8_1181_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_10 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_10) + $signed(sIMD2INT8_1184_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_11 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_11) + $signed(sIMD2INT8_1187_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_12 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_12) + $signed(sIMD2INT8_1190_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_13 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_13) + $signed(sIMD2INT8_1193_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_14 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_14) + $signed(sIMD2INT8_1196_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_15 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_15) + $signed(sIMD2INT8_1199_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_16 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_16) + $signed(sIMD2INT8_1202_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_17 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_17) + $signed(sIMD2INT8_1205_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_18 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_18) + $signed(sIMD2INT8_1208_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_19 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_19) + $signed(sIMD2INT8_1211_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_20 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_20) + $signed(sIMD2INT8_1214_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_21 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_21) + $signed(sIMD2INT8_1217_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_22 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_22) + $signed(sIMD2INT8_1220_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_23 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_23) + $signed(sIMD2INT8_1223_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_24 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_24) + $signed(sIMD2INT8_1226_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_25 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_25) + $signed(sIMD2INT8_1229_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_26 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_26) + $signed(sIMD2INT8_1232_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_27 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_27) + $signed(sIMD2INT8_1235_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_28 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_28) + $signed(sIMD2INT8_1238_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_29 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_29) + $signed(sIMD2INT8_1241_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_30 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_30) + $signed(sIMD2INT8_1244_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_31 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_31) + $signed(sIMD2INT8_1247_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_32 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_32) + $signed(sIMD2INT8_1250_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_33 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_33) + $signed(sIMD2INT8_1253_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_34 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_34) + $signed(sIMD2INT8_1256_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_35 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_35) + $signed(sIMD2INT8_1259_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_36 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_36) + $signed(sIMD2INT8_1262_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_37 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_37) + $signed(sIMD2INT8_1265_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_38 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_38) + $signed(sIMD2INT8_1268_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_39 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_39) + $signed(sIMD2INT8_1271_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_40 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_40) + $signed(sIMD2INT8_1274_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_41 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_41) + $signed(sIMD2INT8_1277_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_42 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_42) + $signed(sIMD2INT8_1280_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_43 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_43) + $signed(sIMD2INT8_1283_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_44 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_44) + $signed(sIMD2INT8_1286_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_45 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_45) + $signed(sIMD2INT8_1289_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_46 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_46) + $signed(sIMD2INT8_1292_ac));
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_pixel_1_47 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_47) + $signed(sIMD2INT8_1295_ac));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_48 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_48) + $signed(tmp_postConv_payload_frame_line_pixel_1_2));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_49 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_49) + $signed(tmp_postConv_payload_frame_line_pixel_1_5));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_50 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_50) + $signed(tmp_postConv_payload_frame_line_pixel_1_8));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_51 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_51) + $signed(tmp_postConv_payload_frame_line_pixel_1_11));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_52 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_52) + $signed(tmp_postConv_payload_frame_line_pixel_1_14));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_53 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_53) + $signed(tmp_postConv_payload_frame_line_pixel_1_17));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_54 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_54) + $signed(tmp_postConv_payload_frame_line_pixel_1_20));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_55 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_55) + $signed(tmp_postConv_payload_frame_line_pixel_1_23));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_56 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_56) + $signed(tmp_postConv_payload_frame_line_pixel_1_26));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_57 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_57) + $signed(tmp_postConv_payload_frame_line_pixel_1_29));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_58 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_58) + $signed(tmp_postConv_payload_frame_line_pixel_1_32));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_59 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_59) + $signed(tmp_postConv_payload_frame_line_pixel_1_35));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_60 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_60) + $signed(tmp_postConv_payload_frame_line_pixel_1_38));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_61 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_61) + $signed(tmp_postConv_payload_frame_line_pixel_1_41));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_62 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_62) + $signed(tmp_postConv_payload_frame_line_pixel_1_44));
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_pixel_1_63 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_63) + $signed(tmp_postConv_payload_frame_line_pixel_1_47));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_64 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_64) + $signed(tmp_postConv_payload_frame_line_pixel_1_50));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_65 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_65) + $signed(tmp_postConv_payload_frame_line_pixel_1_53));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_66 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_66) + $signed(tmp_postConv_payload_frame_line_pixel_1_56));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_67 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_67) + $signed(tmp_postConv_payload_frame_line_pixel_1_59));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_68 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_68) + $signed(tmp_postConv_payload_frame_line_pixel_1_62));
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_pixel_1_69 <= tmp_postConv_payload_frame_line_pixel_1_63;
    end
    if(eventM2sPipes_9_CEs_7) begin
      tmp_postConv_payload_frame_line_pixel_1_70 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_70) + $signed(tmp_postConv_payload_frame_line_pixel_1_66));
    end
    if(eventM2sPipes_9_CEs_7) begin
      tmp_postConv_payload_frame_line_pixel_1_71 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_71) + $signed(tmp_postConv_payload_frame_line_pixel_1_69));
    end
    if(eventM2sPipes_9_CEs_8) begin
      tmp_postConv_payload_frame_line_pixel_1_72 <= ($signed(tmp_tmp_postConv_payload_frame_line_pixel_1_72) + $signed(tmp_tmp_postConv_payload_frame_line_pixel_1_72_1));
    end
    if(eventM2sPipes_9_CEs_0) begin
      tmp_postConv_payload_frame_line_endOfLine <= prevConv_payload_frame_line_endOfLine;
      tmp_postConv_payload_frame_endOfFrame <= prevConv_payload_frame_endOfFrame;
      tmp_postConv_payload_endOfPack <= prevConv_payload_endOfPack;
    end
    if(eventM2sPipes_9_CEs_1) begin
      tmp_postConv_payload_frame_line_endOfLine_1 <= tmp_postConv_payload_frame_line_endOfLine;
      tmp_postConv_payload_frame_endOfFrame_1 <= tmp_postConv_payload_frame_endOfFrame;
      tmp_postConv_payload_endOfPack_1 <= tmp_postConv_payload_endOfPack;
    end
    if(eventM2sPipes_9_CEs_2) begin
      tmp_postConv_payload_frame_line_endOfLine_2 <= tmp_postConv_payload_frame_line_endOfLine_1;
      tmp_postConv_payload_frame_endOfFrame_2 <= tmp_postConv_payload_frame_endOfFrame_1;
      tmp_postConv_payload_endOfPack_2 <= tmp_postConv_payload_endOfPack_1;
    end
    if(eventM2sPipes_9_CEs_3) begin
      tmp_postConv_payload_frame_line_endOfLine_3 <= tmp_postConv_payload_frame_line_endOfLine_2;
      tmp_postConv_payload_frame_endOfFrame_3 <= tmp_postConv_payload_frame_endOfFrame_2;
      tmp_postConv_payload_endOfPack_3 <= tmp_postConv_payload_endOfPack_2;
    end
    if(eventM2sPipes_9_CEs_4) begin
      tmp_postConv_payload_frame_line_endOfLine_4 <= tmp_postConv_payload_frame_line_endOfLine_3;
      tmp_postConv_payload_frame_endOfFrame_4 <= tmp_postConv_payload_frame_endOfFrame_3;
      tmp_postConv_payload_endOfPack_4 <= tmp_postConv_payload_endOfPack_3;
    end
    if(eventM2sPipes_9_CEs_5) begin
      tmp_postConv_payload_frame_line_endOfLine_5 <= tmp_postConv_payload_frame_line_endOfLine_4;
      tmp_postConv_payload_frame_endOfFrame_5 <= tmp_postConv_payload_frame_endOfFrame_4;
      tmp_postConv_payload_endOfPack_5 <= tmp_postConv_payload_endOfPack_4;
    end
    if(eventM2sPipes_9_CEs_6) begin
      tmp_postConv_payload_frame_line_endOfLine_6 <= tmp_postConv_payload_frame_line_endOfLine_5;
      tmp_postConv_payload_frame_endOfFrame_6 <= tmp_postConv_payload_frame_endOfFrame_5;
      tmp_postConv_payload_endOfPack_6 <= tmp_postConv_payload_endOfPack_5;
    end
    if(eventM2sPipes_9_CEs_7) begin
      tmp_postConv_payload_frame_line_endOfLine_7 <= tmp_postConv_payload_frame_line_endOfLine_6;
      tmp_postConv_payload_frame_endOfFrame_7 <= tmp_postConv_payload_frame_endOfFrame_6;
      tmp_postConv_payload_endOfPack_7 <= tmp_postConv_payload_endOfPack_6;
    end
    if(eventM2sPipes_9_CEs_8) begin
      tmp_postConv_payload_frame_line_endOfLine_8 <= tmp_postConv_payload_frame_line_endOfLine_7;
      tmp_postConv_payload_frame_endOfFrame_8 <= tmp_postConv_payload_frame_endOfFrame_7;
      tmp_postConv_payload_endOfPack_8 <= tmp_postConv_payload_endOfPack_7;
    end
    if(postConv_ready) begin
      postConv_rData_frame_line_pixel_0 <= postConv_payload_frame_line_pixel_0;
      postConv_rData_frame_line_pixel_1 <= postConv_payload_frame_line_pixel_1;
      postConv_rData_frame_line_endOfLine <= postConv_payload_frame_line_endOfLine;
      postConv_rData_frame_endOfFrame <= postConv_payload_frame_endOfFrame;
      postConv_rData_endOfPack <= postConv_payload_endOfPack;
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      postConv_rValid <= 1'b0;
    end else begin
      if(postConv_valid) begin
        postConv_rValid <= 1'b1;
      end
      if(postConv_s2mPipe_ready) begin
        postConv_rValid <= 1'b0;
      end
    end
  end


endmodule

module StreamFork_4 (
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_0,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_1,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_2,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_3,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_4,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_5,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_6,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_7,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_8,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_9,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_10,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_11,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_12,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_13,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_14,
  input      [7:0]    io_input_payload_frame_line_pixel_0_0_15,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_0,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_1,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_2,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_3,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_4,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_5,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_6,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_7,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_8,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_9,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_10,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_11,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_12,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_13,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_14,
  input      [7:0]    io_input_payload_frame_line_pixel_0_1_15,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_0,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_1,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_2,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_3,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_4,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_5,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_6,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_7,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_8,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_9,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_10,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_11,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_12,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_13,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_14,
  input      [7:0]    io_input_payload_frame_line_pixel_0_2_15,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_0,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_1,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_2,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_3,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_4,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_5,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_6,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_7,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_8,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_9,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_10,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_11,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_12,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_13,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_14,
  input      [7:0]    io_input_payload_frame_line_pixel_1_0_15,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_0,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_1,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_2,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_3,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_4,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_5,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_6,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_7,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_8,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_9,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_10,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_11,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_12,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_13,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_14,
  input      [7:0]    io_input_payload_frame_line_pixel_1_1_15,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_0,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_1,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_2,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_3,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_4,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_5,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_6,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_7,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_8,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_9,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_10,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_11,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_12,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_13,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_14,
  input      [7:0]    io_input_payload_frame_line_pixel_1_2_15,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_0,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_1,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_2,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_3,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_4,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_5,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_6,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_7,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_8,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_9,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_10,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_11,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_12,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_13,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_14,
  input      [7:0]    io_input_payload_frame_line_pixel_2_0_15,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_0,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_1,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_2,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_3,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_4,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_5,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_6,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_7,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_8,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_9,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_10,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_11,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_12,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_13,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_14,
  input      [7:0]    io_input_payload_frame_line_pixel_2_1_15,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_0,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_1,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_2,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_3,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_4,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_5,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_6,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_7,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_8,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_9,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_10,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_11,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_12,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_13,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_14,
  input      [7:0]    io_input_payload_frame_line_pixel_2_2_15,
  input               io_input_payload_frame_line_endOfLine,
  input               io_input_payload_frame_endOfFrame,
  input               io_input_payload_endOfPack,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2_2_15,
  output              io_outputs_0_payload_frame_line_endOfLine,
  output              io_outputs_0_payload_frame_endOfFrame,
  output              io_outputs_0_payload_endOfPack,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2_2_15,
  output              io_outputs_1_payload_frame_line_endOfLine,
  output              io_outputs_1_payload_frame_endOfFrame,
  output              io_outputs_1_payload_endOfPack,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_2_payload_frame_line_pixel_2_2_15,
  output              io_outputs_2_payload_frame_line_endOfLine,
  output              io_outputs_2_payload_frame_endOfFrame,
  output              io_outputs_2_payload_endOfPack,
  output              io_outputs_3_valid,
  input               io_outputs_3_ready,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_3_payload_frame_line_pixel_2_2_15,
  output              io_outputs_3_payload_frame_line_endOfLine,
  output              io_outputs_3_payload_frame_endOfFrame,
  output              io_outputs_3_payload_endOfPack,
  output              io_outputs_4_valid,
  input               io_outputs_4_ready,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_4_payload_frame_line_pixel_2_2_15,
  output              io_outputs_4_payload_frame_line_endOfLine,
  output              io_outputs_4_payload_frame_endOfFrame,
  output              io_outputs_4_payload_endOfPack,
  output              io_outputs_5_valid,
  input               io_outputs_5_ready,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_5_payload_frame_line_pixel_2_2_15,
  output              io_outputs_5_payload_frame_line_endOfLine,
  output              io_outputs_5_payload_frame_endOfFrame,
  output              io_outputs_5_payload_endOfPack,
  output              io_outputs_6_valid,
  input               io_outputs_6_ready,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_6_payload_frame_line_pixel_2_2_15,
  output              io_outputs_6_payload_frame_line_endOfLine,
  output              io_outputs_6_payload_frame_endOfFrame,
  output              io_outputs_6_payload_endOfPack,
  output              io_outputs_7_valid,
  input               io_outputs_7_ready,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_0_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_1_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_0_2_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_0_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_1_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_1_2_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_0_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_1_15,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_0,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_1,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_2,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_3,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_4,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_5,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_6,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_7,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_8,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_9,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_10,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_11,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_12,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_13,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_14,
  output     [7:0]    io_outputs_7_payload_frame_line_pixel_2_2_15,
  output              io_outputs_7_payload_frame_line_endOfLine,
  output              io_outputs_7_payload_frame_endOfFrame,
  output              io_outputs_7_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 tmp_io_outputs_0_valid;
  reg                 tmp_io_outputs_1_valid;
  reg                 tmp_io_outputs_2_valid;
  reg                 tmp_io_outputs_3_valid;
  reg                 tmp_io_outputs_4_valid;
  reg                 tmp_io_outputs_5_valid;
  reg                 tmp_io_outputs_6_valid;
  reg                 tmp_io_outputs_7_valid;
  wire                when_Stream_l825;
  wire                when_Stream_l825_1;
  wire                when_Stream_l825_2;
  wire                when_Stream_l825_3;
  wire                when_Stream_l825_4;
  wire                when_Stream_l825_5;
  wire                when_Stream_l825_6;
  wire                when_Stream_l825_7;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;
  wire                io_outputs_2_fire;
  wire                io_outputs_3_fire;
  wire                io_outputs_4_fire;
  wire                io_outputs_5_fire;
  wire                io_outputs_6_fire;
  wire                io_outputs_7_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l825) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_1) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_2) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_3) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_4) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_5) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_6) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_7) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l825 = ((! io_outputs_0_ready) && tmp_io_outputs_0_valid);
  assign when_Stream_l825_1 = ((! io_outputs_1_ready) && tmp_io_outputs_1_valid);
  assign when_Stream_l825_2 = ((! io_outputs_2_ready) && tmp_io_outputs_2_valid);
  assign when_Stream_l825_3 = ((! io_outputs_3_ready) && tmp_io_outputs_3_valid);
  assign when_Stream_l825_4 = ((! io_outputs_4_ready) && tmp_io_outputs_4_valid);
  assign when_Stream_l825_5 = ((! io_outputs_5_ready) && tmp_io_outputs_5_valid);
  assign when_Stream_l825_6 = ((! io_outputs_6_ready) && tmp_io_outputs_6_valid);
  assign when_Stream_l825_7 = ((! io_outputs_7_ready) && tmp_io_outputs_7_valid);
  assign io_outputs_0_valid = (io_input_valid && tmp_io_outputs_0_valid);
  assign io_outputs_0_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_0_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_0_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_0_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_0_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_0_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_0_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_0_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_0_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_0_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_0_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_0_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_0_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_0_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_0_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_0_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_0_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_0_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_0_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_0_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_0_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_0_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_0_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_0_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_0_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_0_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_0_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_0_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_0_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_0_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_0_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_0_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_0_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_0_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_0_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_0_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_0_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_0_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_0_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_0_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_0_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_0_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_0_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_0_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_0_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_0_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_0_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_0_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_0_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_0_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_0_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_0_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_0_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_0_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_0_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_0_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_0_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_0_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_0_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_0_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_0_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_0_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_0_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_0_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_0_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_0_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_0_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_0_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_0_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_0_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_0_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_0_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_0_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_0_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_0_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_0_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_0_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_0_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_0_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_0_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_0_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_0_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_0_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_0_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_0_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_0_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_0_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_0_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_0_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_0_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_0_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_0_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_0_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_0_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_0_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_0_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_0_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_0_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_0_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_0_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_0_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_0_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_0_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_0_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_0_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_0_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_0_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_0_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_0_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_0_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_0_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_0_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_0_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_0_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_0_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_0_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_0_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_0_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_0_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_0_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_0_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_0_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_0_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_0_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_0_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_0_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_0_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_0_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_0_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_0_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_0_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_0_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_0_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_0_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_0_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_0_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_0_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_0_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_0_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_0_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_0_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_0_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_0_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_0_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_0_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_0_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_0_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && tmp_io_outputs_1_valid);
  assign io_outputs_1_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_1_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_1_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_1_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_1_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_1_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_1_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_1_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_1_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_1_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_1_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_1_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_1_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_1_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_1_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_1_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_1_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_1_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_1_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_1_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_1_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_1_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_1_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_1_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_1_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_1_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_1_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_1_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_1_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_1_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_1_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_1_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_1_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_1_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_1_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_1_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_1_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_1_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_1_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_1_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_1_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_1_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_1_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_1_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_1_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_1_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_1_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_1_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_1_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_1_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_1_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_1_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_1_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_1_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_1_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_1_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_1_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_1_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_1_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_1_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_1_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_1_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_1_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_1_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_1_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_1_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_1_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_1_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_1_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_1_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_1_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_1_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_1_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_1_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_1_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_1_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_1_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_1_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_1_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_1_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_1_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_1_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_1_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_1_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_1_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_1_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_1_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_1_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_1_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_1_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_1_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_1_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_1_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_1_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_1_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_1_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_1_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_1_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_1_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_1_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_1_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_1_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_1_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_1_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_1_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_1_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_1_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_1_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_1_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_1_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_1_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_1_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_1_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_1_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_1_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_1_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_1_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_1_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_1_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_1_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_1_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_1_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_1_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_1_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_1_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_1_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_1_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_1_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_1_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_1_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_1_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_1_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_1_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_1_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_1_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_1_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_1_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_1_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_1_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_1_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_1_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_1_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_1_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_1_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_1_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_1_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_1_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  assign io_outputs_2_valid = (io_input_valid && tmp_io_outputs_2_valid);
  assign io_outputs_2_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_2_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_2_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_2_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_2_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_2_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_2_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_2_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_2_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_2_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_2_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_2_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_2_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_2_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_2_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_2_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_2_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_2_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_2_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_2_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_2_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_2_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_2_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_2_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_2_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_2_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_2_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_2_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_2_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_2_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_2_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_2_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_2_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_2_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_2_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_2_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_2_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_2_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_2_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_2_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_2_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_2_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_2_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_2_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_2_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_2_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_2_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_2_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_2_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_2_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_2_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_2_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_2_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_2_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_2_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_2_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_2_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_2_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_2_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_2_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_2_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_2_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_2_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_2_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_2_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_2_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_2_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_2_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_2_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_2_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_2_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_2_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_2_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_2_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_2_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_2_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_2_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_2_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_2_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_2_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_2_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_2_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_2_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_2_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_2_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_2_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_2_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_2_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_2_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_2_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_2_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_2_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_2_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_2_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_2_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_2_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_2_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_2_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_2_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_2_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_2_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_2_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_2_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_2_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_2_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_2_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_2_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_2_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_2_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_2_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_2_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_2_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_2_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_2_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_2_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_2_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_2_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_2_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_2_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_2_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_2_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_2_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_2_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_2_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_2_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_2_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_2_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_2_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_2_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_2_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_2_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_2_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_2_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_2_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_2_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_2_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_2_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_2_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_2_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_2_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_2_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_2_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_2_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_2_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_2_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_2_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_2_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_2_fire = (io_outputs_2_valid && io_outputs_2_ready);
  assign io_outputs_3_valid = (io_input_valid && tmp_io_outputs_3_valid);
  assign io_outputs_3_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_3_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_3_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_3_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_3_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_3_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_3_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_3_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_3_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_3_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_3_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_3_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_3_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_3_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_3_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_3_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_3_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_3_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_3_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_3_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_3_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_3_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_3_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_3_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_3_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_3_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_3_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_3_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_3_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_3_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_3_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_3_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_3_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_3_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_3_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_3_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_3_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_3_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_3_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_3_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_3_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_3_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_3_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_3_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_3_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_3_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_3_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_3_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_3_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_3_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_3_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_3_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_3_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_3_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_3_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_3_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_3_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_3_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_3_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_3_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_3_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_3_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_3_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_3_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_3_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_3_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_3_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_3_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_3_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_3_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_3_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_3_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_3_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_3_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_3_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_3_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_3_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_3_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_3_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_3_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_3_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_3_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_3_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_3_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_3_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_3_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_3_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_3_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_3_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_3_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_3_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_3_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_3_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_3_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_3_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_3_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_3_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_3_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_3_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_3_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_3_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_3_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_3_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_3_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_3_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_3_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_3_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_3_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_3_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_3_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_3_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_3_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_3_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_3_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_3_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_3_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_3_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_3_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_3_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_3_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_3_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_3_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_3_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_3_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_3_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_3_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_3_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_3_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_3_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_3_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_3_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_3_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_3_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_3_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_3_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_3_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_3_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_3_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_3_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_3_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_3_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_3_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_3_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_3_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_3_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_3_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_3_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_3_fire = (io_outputs_3_valid && io_outputs_3_ready);
  assign io_outputs_4_valid = (io_input_valid && tmp_io_outputs_4_valid);
  assign io_outputs_4_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_4_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_4_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_4_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_4_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_4_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_4_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_4_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_4_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_4_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_4_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_4_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_4_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_4_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_4_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_4_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_4_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_4_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_4_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_4_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_4_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_4_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_4_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_4_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_4_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_4_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_4_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_4_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_4_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_4_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_4_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_4_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_4_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_4_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_4_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_4_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_4_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_4_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_4_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_4_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_4_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_4_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_4_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_4_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_4_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_4_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_4_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_4_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_4_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_4_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_4_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_4_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_4_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_4_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_4_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_4_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_4_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_4_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_4_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_4_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_4_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_4_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_4_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_4_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_4_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_4_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_4_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_4_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_4_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_4_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_4_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_4_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_4_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_4_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_4_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_4_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_4_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_4_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_4_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_4_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_4_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_4_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_4_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_4_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_4_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_4_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_4_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_4_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_4_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_4_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_4_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_4_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_4_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_4_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_4_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_4_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_4_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_4_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_4_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_4_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_4_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_4_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_4_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_4_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_4_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_4_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_4_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_4_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_4_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_4_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_4_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_4_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_4_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_4_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_4_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_4_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_4_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_4_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_4_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_4_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_4_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_4_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_4_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_4_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_4_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_4_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_4_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_4_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_4_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_4_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_4_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_4_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_4_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_4_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_4_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_4_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_4_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_4_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_4_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_4_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_4_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_4_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_4_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_4_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_4_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_4_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_4_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_4_fire = (io_outputs_4_valid && io_outputs_4_ready);
  assign io_outputs_5_valid = (io_input_valid && tmp_io_outputs_5_valid);
  assign io_outputs_5_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_5_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_5_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_5_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_5_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_5_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_5_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_5_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_5_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_5_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_5_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_5_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_5_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_5_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_5_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_5_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_5_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_5_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_5_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_5_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_5_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_5_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_5_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_5_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_5_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_5_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_5_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_5_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_5_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_5_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_5_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_5_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_5_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_5_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_5_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_5_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_5_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_5_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_5_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_5_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_5_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_5_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_5_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_5_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_5_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_5_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_5_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_5_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_5_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_5_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_5_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_5_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_5_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_5_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_5_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_5_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_5_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_5_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_5_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_5_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_5_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_5_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_5_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_5_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_5_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_5_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_5_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_5_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_5_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_5_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_5_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_5_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_5_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_5_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_5_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_5_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_5_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_5_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_5_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_5_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_5_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_5_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_5_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_5_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_5_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_5_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_5_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_5_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_5_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_5_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_5_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_5_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_5_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_5_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_5_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_5_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_5_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_5_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_5_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_5_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_5_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_5_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_5_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_5_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_5_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_5_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_5_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_5_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_5_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_5_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_5_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_5_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_5_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_5_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_5_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_5_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_5_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_5_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_5_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_5_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_5_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_5_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_5_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_5_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_5_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_5_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_5_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_5_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_5_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_5_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_5_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_5_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_5_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_5_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_5_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_5_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_5_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_5_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_5_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_5_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_5_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_5_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_5_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_5_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_5_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_5_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_5_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_5_fire = (io_outputs_5_valid && io_outputs_5_ready);
  assign io_outputs_6_valid = (io_input_valid && tmp_io_outputs_6_valid);
  assign io_outputs_6_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_6_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_6_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_6_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_6_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_6_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_6_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_6_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_6_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_6_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_6_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_6_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_6_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_6_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_6_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_6_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_6_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_6_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_6_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_6_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_6_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_6_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_6_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_6_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_6_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_6_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_6_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_6_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_6_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_6_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_6_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_6_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_6_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_6_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_6_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_6_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_6_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_6_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_6_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_6_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_6_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_6_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_6_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_6_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_6_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_6_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_6_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_6_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_6_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_6_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_6_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_6_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_6_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_6_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_6_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_6_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_6_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_6_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_6_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_6_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_6_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_6_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_6_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_6_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_6_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_6_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_6_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_6_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_6_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_6_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_6_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_6_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_6_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_6_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_6_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_6_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_6_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_6_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_6_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_6_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_6_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_6_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_6_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_6_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_6_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_6_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_6_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_6_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_6_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_6_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_6_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_6_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_6_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_6_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_6_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_6_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_6_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_6_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_6_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_6_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_6_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_6_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_6_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_6_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_6_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_6_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_6_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_6_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_6_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_6_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_6_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_6_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_6_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_6_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_6_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_6_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_6_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_6_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_6_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_6_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_6_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_6_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_6_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_6_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_6_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_6_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_6_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_6_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_6_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_6_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_6_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_6_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_6_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_6_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_6_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_6_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_6_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_6_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_6_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_6_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_6_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_6_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_6_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_6_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_6_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_6_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_6_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_6_fire = (io_outputs_6_valid && io_outputs_6_ready);
  assign io_outputs_7_valid = (io_input_valid && tmp_io_outputs_7_valid);
  assign io_outputs_7_payload_frame_line_pixel_0_0_0 = io_input_payload_frame_line_pixel_0_0_0;
  assign io_outputs_7_payload_frame_line_pixel_0_0_1 = io_input_payload_frame_line_pixel_0_0_1;
  assign io_outputs_7_payload_frame_line_pixel_0_0_2 = io_input_payload_frame_line_pixel_0_0_2;
  assign io_outputs_7_payload_frame_line_pixel_0_0_3 = io_input_payload_frame_line_pixel_0_0_3;
  assign io_outputs_7_payload_frame_line_pixel_0_0_4 = io_input_payload_frame_line_pixel_0_0_4;
  assign io_outputs_7_payload_frame_line_pixel_0_0_5 = io_input_payload_frame_line_pixel_0_0_5;
  assign io_outputs_7_payload_frame_line_pixel_0_0_6 = io_input_payload_frame_line_pixel_0_0_6;
  assign io_outputs_7_payload_frame_line_pixel_0_0_7 = io_input_payload_frame_line_pixel_0_0_7;
  assign io_outputs_7_payload_frame_line_pixel_0_0_8 = io_input_payload_frame_line_pixel_0_0_8;
  assign io_outputs_7_payload_frame_line_pixel_0_0_9 = io_input_payload_frame_line_pixel_0_0_9;
  assign io_outputs_7_payload_frame_line_pixel_0_0_10 = io_input_payload_frame_line_pixel_0_0_10;
  assign io_outputs_7_payload_frame_line_pixel_0_0_11 = io_input_payload_frame_line_pixel_0_0_11;
  assign io_outputs_7_payload_frame_line_pixel_0_0_12 = io_input_payload_frame_line_pixel_0_0_12;
  assign io_outputs_7_payload_frame_line_pixel_0_0_13 = io_input_payload_frame_line_pixel_0_0_13;
  assign io_outputs_7_payload_frame_line_pixel_0_0_14 = io_input_payload_frame_line_pixel_0_0_14;
  assign io_outputs_7_payload_frame_line_pixel_0_0_15 = io_input_payload_frame_line_pixel_0_0_15;
  assign io_outputs_7_payload_frame_line_pixel_0_1_0 = io_input_payload_frame_line_pixel_0_1_0;
  assign io_outputs_7_payload_frame_line_pixel_0_1_1 = io_input_payload_frame_line_pixel_0_1_1;
  assign io_outputs_7_payload_frame_line_pixel_0_1_2 = io_input_payload_frame_line_pixel_0_1_2;
  assign io_outputs_7_payload_frame_line_pixel_0_1_3 = io_input_payload_frame_line_pixel_0_1_3;
  assign io_outputs_7_payload_frame_line_pixel_0_1_4 = io_input_payload_frame_line_pixel_0_1_4;
  assign io_outputs_7_payload_frame_line_pixel_0_1_5 = io_input_payload_frame_line_pixel_0_1_5;
  assign io_outputs_7_payload_frame_line_pixel_0_1_6 = io_input_payload_frame_line_pixel_0_1_6;
  assign io_outputs_7_payload_frame_line_pixel_0_1_7 = io_input_payload_frame_line_pixel_0_1_7;
  assign io_outputs_7_payload_frame_line_pixel_0_1_8 = io_input_payload_frame_line_pixel_0_1_8;
  assign io_outputs_7_payload_frame_line_pixel_0_1_9 = io_input_payload_frame_line_pixel_0_1_9;
  assign io_outputs_7_payload_frame_line_pixel_0_1_10 = io_input_payload_frame_line_pixel_0_1_10;
  assign io_outputs_7_payload_frame_line_pixel_0_1_11 = io_input_payload_frame_line_pixel_0_1_11;
  assign io_outputs_7_payload_frame_line_pixel_0_1_12 = io_input_payload_frame_line_pixel_0_1_12;
  assign io_outputs_7_payload_frame_line_pixel_0_1_13 = io_input_payload_frame_line_pixel_0_1_13;
  assign io_outputs_7_payload_frame_line_pixel_0_1_14 = io_input_payload_frame_line_pixel_0_1_14;
  assign io_outputs_7_payload_frame_line_pixel_0_1_15 = io_input_payload_frame_line_pixel_0_1_15;
  assign io_outputs_7_payload_frame_line_pixel_0_2_0 = io_input_payload_frame_line_pixel_0_2_0;
  assign io_outputs_7_payload_frame_line_pixel_0_2_1 = io_input_payload_frame_line_pixel_0_2_1;
  assign io_outputs_7_payload_frame_line_pixel_0_2_2 = io_input_payload_frame_line_pixel_0_2_2;
  assign io_outputs_7_payload_frame_line_pixel_0_2_3 = io_input_payload_frame_line_pixel_0_2_3;
  assign io_outputs_7_payload_frame_line_pixel_0_2_4 = io_input_payload_frame_line_pixel_0_2_4;
  assign io_outputs_7_payload_frame_line_pixel_0_2_5 = io_input_payload_frame_line_pixel_0_2_5;
  assign io_outputs_7_payload_frame_line_pixel_0_2_6 = io_input_payload_frame_line_pixel_0_2_6;
  assign io_outputs_7_payload_frame_line_pixel_0_2_7 = io_input_payload_frame_line_pixel_0_2_7;
  assign io_outputs_7_payload_frame_line_pixel_0_2_8 = io_input_payload_frame_line_pixel_0_2_8;
  assign io_outputs_7_payload_frame_line_pixel_0_2_9 = io_input_payload_frame_line_pixel_0_2_9;
  assign io_outputs_7_payload_frame_line_pixel_0_2_10 = io_input_payload_frame_line_pixel_0_2_10;
  assign io_outputs_7_payload_frame_line_pixel_0_2_11 = io_input_payload_frame_line_pixel_0_2_11;
  assign io_outputs_7_payload_frame_line_pixel_0_2_12 = io_input_payload_frame_line_pixel_0_2_12;
  assign io_outputs_7_payload_frame_line_pixel_0_2_13 = io_input_payload_frame_line_pixel_0_2_13;
  assign io_outputs_7_payload_frame_line_pixel_0_2_14 = io_input_payload_frame_line_pixel_0_2_14;
  assign io_outputs_7_payload_frame_line_pixel_0_2_15 = io_input_payload_frame_line_pixel_0_2_15;
  assign io_outputs_7_payload_frame_line_pixel_1_0_0 = io_input_payload_frame_line_pixel_1_0_0;
  assign io_outputs_7_payload_frame_line_pixel_1_0_1 = io_input_payload_frame_line_pixel_1_0_1;
  assign io_outputs_7_payload_frame_line_pixel_1_0_2 = io_input_payload_frame_line_pixel_1_0_2;
  assign io_outputs_7_payload_frame_line_pixel_1_0_3 = io_input_payload_frame_line_pixel_1_0_3;
  assign io_outputs_7_payload_frame_line_pixel_1_0_4 = io_input_payload_frame_line_pixel_1_0_4;
  assign io_outputs_7_payload_frame_line_pixel_1_0_5 = io_input_payload_frame_line_pixel_1_0_5;
  assign io_outputs_7_payload_frame_line_pixel_1_0_6 = io_input_payload_frame_line_pixel_1_0_6;
  assign io_outputs_7_payload_frame_line_pixel_1_0_7 = io_input_payload_frame_line_pixel_1_0_7;
  assign io_outputs_7_payload_frame_line_pixel_1_0_8 = io_input_payload_frame_line_pixel_1_0_8;
  assign io_outputs_7_payload_frame_line_pixel_1_0_9 = io_input_payload_frame_line_pixel_1_0_9;
  assign io_outputs_7_payload_frame_line_pixel_1_0_10 = io_input_payload_frame_line_pixel_1_0_10;
  assign io_outputs_7_payload_frame_line_pixel_1_0_11 = io_input_payload_frame_line_pixel_1_0_11;
  assign io_outputs_7_payload_frame_line_pixel_1_0_12 = io_input_payload_frame_line_pixel_1_0_12;
  assign io_outputs_7_payload_frame_line_pixel_1_0_13 = io_input_payload_frame_line_pixel_1_0_13;
  assign io_outputs_7_payload_frame_line_pixel_1_0_14 = io_input_payload_frame_line_pixel_1_0_14;
  assign io_outputs_7_payload_frame_line_pixel_1_0_15 = io_input_payload_frame_line_pixel_1_0_15;
  assign io_outputs_7_payload_frame_line_pixel_1_1_0 = io_input_payload_frame_line_pixel_1_1_0;
  assign io_outputs_7_payload_frame_line_pixel_1_1_1 = io_input_payload_frame_line_pixel_1_1_1;
  assign io_outputs_7_payload_frame_line_pixel_1_1_2 = io_input_payload_frame_line_pixel_1_1_2;
  assign io_outputs_7_payload_frame_line_pixel_1_1_3 = io_input_payload_frame_line_pixel_1_1_3;
  assign io_outputs_7_payload_frame_line_pixel_1_1_4 = io_input_payload_frame_line_pixel_1_1_4;
  assign io_outputs_7_payload_frame_line_pixel_1_1_5 = io_input_payload_frame_line_pixel_1_1_5;
  assign io_outputs_7_payload_frame_line_pixel_1_1_6 = io_input_payload_frame_line_pixel_1_1_6;
  assign io_outputs_7_payload_frame_line_pixel_1_1_7 = io_input_payload_frame_line_pixel_1_1_7;
  assign io_outputs_7_payload_frame_line_pixel_1_1_8 = io_input_payload_frame_line_pixel_1_1_8;
  assign io_outputs_7_payload_frame_line_pixel_1_1_9 = io_input_payload_frame_line_pixel_1_1_9;
  assign io_outputs_7_payload_frame_line_pixel_1_1_10 = io_input_payload_frame_line_pixel_1_1_10;
  assign io_outputs_7_payload_frame_line_pixel_1_1_11 = io_input_payload_frame_line_pixel_1_1_11;
  assign io_outputs_7_payload_frame_line_pixel_1_1_12 = io_input_payload_frame_line_pixel_1_1_12;
  assign io_outputs_7_payload_frame_line_pixel_1_1_13 = io_input_payload_frame_line_pixel_1_1_13;
  assign io_outputs_7_payload_frame_line_pixel_1_1_14 = io_input_payload_frame_line_pixel_1_1_14;
  assign io_outputs_7_payload_frame_line_pixel_1_1_15 = io_input_payload_frame_line_pixel_1_1_15;
  assign io_outputs_7_payload_frame_line_pixel_1_2_0 = io_input_payload_frame_line_pixel_1_2_0;
  assign io_outputs_7_payload_frame_line_pixel_1_2_1 = io_input_payload_frame_line_pixel_1_2_1;
  assign io_outputs_7_payload_frame_line_pixel_1_2_2 = io_input_payload_frame_line_pixel_1_2_2;
  assign io_outputs_7_payload_frame_line_pixel_1_2_3 = io_input_payload_frame_line_pixel_1_2_3;
  assign io_outputs_7_payload_frame_line_pixel_1_2_4 = io_input_payload_frame_line_pixel_1_2_4;
  assign io_outputs_7_payload_frame_line_pixel_1_2_5 = io_input_payload_frame_line_pixel_1_2_5;
  assign io_outputs_7_payload_frame_line_pixel_1_2_6 = io_input_payload_frame_line_pixel_1_2_6;
  assign io_outputs_7_payload_frame_line_pixel_1_2_7 = io_input_payload_frame_line_pixel_1_2_7;
  assign io_outputs_7_payload_frame_line_pixel_1_2_8 = io_input_payload_frame_line_pixel_1_2_8;
  assign io_outputs_7_payload_frame_line_pixel_1_2_9 = io_input_payload_frame_line_pixel_1_2_9;
  assign io_outputs_7_payload_frame_line_pixel_1_2_10 = io_input_payload_frame_line_pixel_1_2_10;
  assign io_outputs_7_payload_frame_line_pixel_1_2_11 = io_input_payload_frame_line_pixel_1_2_11;
  assign io_outputs_7_payload_frame_line_pixel_1_2_12 = io_input_payload_frame_line_pixel_1_2_12;
  assign io_outputs_7_payload_frame_line_pixel_1_2_13 = io_input_payload_frame_line_pixel_1_2_13;
  assign io_outputs_7_payload_frame_line_pixel_1_2_14 = io_input_payload_frame_line_pixel_1_2_14;
  assign io_outputs_7_payload_frame_line_pixel_1_2_15 = io_input_payload_frame_line_pixel_1_2_15;
  assign io_outputs_7_payload_frame_line_pixel_2_0_0 = io_input_payload_frame_line_pixel_2_0_0;
  assign io_outputs_7_payload_frame_line_pixel_2_0_1 = io_input_payload_frame_line_pixel_2_0_1;
  assign io_outputs_7_payload_frame_line_pixel_2_0_2 = io_input_payload_frame_line_pixel_2_0_2;
  assign io_outputs_7_payload_frame_line_pixel_2_0_3 = io_input_payload_frame_line_pixel_2_0_3;
  assign io_outputs_7_payload_frame_line_pixel_2_0_4 = io_input_payload_frame_line_pixel_2_0_4;
  assign io_outputs_7_payload_frame_line_pixel_2_0_5 = io_input_payload_frame_line_pixel_2_0_5;
  assign io_outputs_7_payload_frame_line_pixel_2_0_6 = io_input_payload_frame_line_pixel_2_0_6;
  assign io_outputs_7_payload_frame_line_pixel_2_0_7 = io_input_payload_frame_line_pixel_2_0_7;
  assign io_outputs_7_payload_frame_line_pixel_2_0_8 = io_input_payload_frame_line_pixel_2_0_8;
  assign io_outputs_7_payload_frame_line_pixel_2_0_9 = io_input_payload_frame_line_pixel_2_0_9;
  assign io_outputs_7_payload_frame_line_pixel_2_0_10 = io_input_payload_frame_line_pixel_2_0_10;
  assign io_outputs_7_payload_frame_line_pixel_2_0_11 = io_input_payload_frame_line_pixel_2_0_11;
  assign io_outputs_7_payload_frame_line_pixel_2_0_12 = io_input_payload_frame_line_pixel_2_0_12;
  assign io_outputs_7_payload_frame_line_pixel_2_0_13 = io_input_payload_frame_line_pixel_2_0_13;
  assign io_outputs_7_payload_frame_line_pixel_2_0_14 = io_input_payload_frame_line_pixel_2_0_14;
  assign io_outputs_7_payload_frame_line_pixel_2_0_15 = io_input_payload_frame_line_pixel_2_0_15;
  assign io_outputs_7_payload_frame_line_pixel_2_1_0 = io_input_payload_frame_line_pixel_2_1_0;
  assign io_outputs_7_payload_frame_line_pixel_2_1_1 = io_input_payload_frame_line_pixel_2_1_1;
  assign io_outputs_7_payload_frame_line_pixel_2_1_2 = io_input_payload_frame_line_pixel_2_1_2;
  assign io_outputs_7_payload_frame_line_pixel_2_1_3 = io_input_payload_frame_line_pixel_2_1_3;
  assign io_outputs_7_payload_frame_line_pixel_2_1_4 = io_input_payload_frame_line_pixel_2_1_4;
  assign io_outputs_7_payload_frame_line_pixel_2_1_5 = io_input_payload_frame_line_pixel_2_1_5;
  assign io_outputs_7_payload_frame_line_pixel_2_1_6 = io_input_payload_frame_line_pixel_2_1_6;
  assign io_outputs_7_payload_frame_line_pixel_2_1_7 = io_input_payload_frame_line_pixel_2_1_7;
  assign io_outputs_7_payload_frame_line_pixel_2_1_8 = io_input_payload_frame_line_pixel_2_1_8;
  assign io_outputs_7_payload_frame_line_pixel_2_1_9 = io_input_payload_frame_line_pixel_2_1_9;
  assign io_outputs_7_payload_frame_line_pixel_2_1_10 = io_input_payload_frame_line_pixel_2_1_10;
  assign io_outputs_7_payload_frame_line_pixel_2_1_11 = io_input_payload_frame_line_pixel_2_1_11;
  assign io_outputs_7_payload_frame_line_pixel_2_1_12 = io_input_payload_frame_line_pixel_2_1_12;
  assign io_outputs_7_payload_frame_line_pixel_2_1_13 = io_input_payload_frame_line_pixel_2_1_13;
  assign io_outputs_7_payload_frame_line_pixel_2_1_14 = io_input_payload_frame_line_pixel_2_1_14;
  assign io_outputs_7_payload_frame_line_pixel_2_1_15 = io_input_payload_frame_line_pixel_2_1_15;
  assign io_outputs_7_payload_frame_line_pixel_2_2_0 = io_input_payload_frame_line_pixel_2_2_0;
  assign io_outputs_7_payload_frame_line_pixel_2_2_1 = io_input_payload_frame_line_pixel_2_2_1;
  assign io_outputs_7_payload_frame_line_pixel_2_2_2 = io_input_payload_frame_line_pixel_2_2_2;
  assign io_outputs_7_payload_frame_line_pixel_2_2_3 = io_input_payload_frame_line_pixel_2_2_3;
  assign io_outputs_7_payload_frame_line_pixel_2_2_4 = io_input_payload_frame_line_pixel_2_2_4;
  assign io_outputs_7_payload_frame_line_pixel_2_2_5 = io_input_payload_frame_line_pixel_2_2_5;
  assign io_outputs_7_payload_frame_line_pixel_2_2_6 = io_input_payload_frame_line_pixel_2_2_6;
  assign io_outputs_7_payload_frame_line_pixel_2_2_7 = io_input_payload_frame_line_pixel_2_2_7;
  assign io_outputs_7_payload_frame_line_pixel_2_2_8 = io_input_payload_frame_line_pixel_2_2_8;
  assign io_outputs_7_payload_frame_line_pixel_2_2_9 = io_input_payload_frame_line_pixel_2_2_9;
  assign io_outputs_7_payload_frame_line_pixel_2_2_10 = io_input_payload_frame_line_pixel_2_2_10;
  assign io_outputs_7_payload_frame_line_pixel_2_2_11 = io_input_payload_frame_line_pixel_2_2_11;
  assign io_outputs_7_payload_frame_line_pixel_2_2_12 = io_input_payload_frame_line_pixel_2_2_12;
  assign io_outputs_7_payload_frame_line_pixel_2_2_13 = io_input_payload_frame_line_pixel_2_2_13;
  assign io_outputs_7_payload_frame_line_pixel_2_2_14 = io_input_payload_frame_line_pixel_2_2_14;
  assign io_outputs_7_payload_frame_line_pixel_2_2_15 = io_input_payload_frame_line_pixel_2_2_15;
  assign io_outputs_7_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_7_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_7_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_7_fire = (io_outputs_7_valid && io_outputs_7_ready);
  always @(posedge clk) begin
    if(reset) begin
      tmp_io_outputs_0_valid <= 1'b1;
      tmp_io_outputs_1_valid <= 1'b1;
      tmp_io_outputs_2_valid <= 1'b1;
      tmp_io_outputs_3_valid <= 1'b1;
      tmp_io_outputs_4_valid <= 1'b1;
      tmp_io_outputs_5_valid <= 1'b1;
      tmp_io_outputs_6_valid <= 1'b1;
      tmp_io_outputs_7_valid <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        tmp_io_outputs_0_valid <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        tmp_io_outputs_1_valid <= 1'b0;
      end
      if(io_outputs_2_fire) begin
        tmp_io_outputs_2_valid <= 1'b0;
      end
      if(io_outputs_3_fire) begin
        tmp_io_outputs_3_valid <= 1'b0;
      end
      if(io_outputs_4_fire) begin
        tmp_io_outputs_4_valid <= 1'b0;
      end
      if(io_outputs_5_fire) begin
        tmp_io_outputs_5_valid <= 1'b0;
      end
      if(io_outputs_6_fire) begin
        tmp_io_outputs_6_valid <= 1'b0;
      end
      if(io_outputs_7_fire) begin
        tmp_io_outputs_7_valid <= 1'b0;
      end
      if(io_input_ready) begin
        tmp_io_outputs_0_valid <= 1'b1;
        tmp_io_outputs_1_valid <= 1'b1;
        tmp_io_outputs_2_valid <= 1'b1;
        tmp_io_outputs_3_valid <= 1'b1;
        tmp_io_outputs_4_valid <= 1'b1;
        tmp_io_outputs_5_valid <= 1'b1;
        tmp_io_outputs_6_valid <= 1'b1;
        tmp_io_outputs_7_valid <= 1'b1;
      end
    end
  end


endmodule

module SlidingWindowSame (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 line_videoOut_ready;
  reg                 pixel_videoOut_ready;
  wire                line_videoIn_ready;
  wire                line_videoOut_valid;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_0;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_1;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_2;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_3;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_4;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_5;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_6;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_7;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_8;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_9;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_10;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_11;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_12;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_13;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_14;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_15;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_0;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_1;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_2;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_3;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_4;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_5;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_6;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_7;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_8;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_9;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_10;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_11;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_12;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_13;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_14;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_15;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_0;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_1;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_2;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_3;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_4;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_5;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_6;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_7;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_8;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_9;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_10;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_11;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_12;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_13;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_14;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_2_15;
  wire                line_videoOut_payload_frame_line_endOfLine;
  wire                line_videoOut_payload_frame_endOfFrame;
  wire                line_videoOut_payload_endOfPack;
  wire                pixel_videoIn_ready;
  wire                pixel_videoOut_valid;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_2_2_15;
  wire                pixel_videoOut_payload_frame_line_endOfLine;
  wire                pixel_videoOut_payload_frame_endOfFrame;
  wire                pixel_videoOut_payload_endOfPack;
  wire                pixelOut_valid;
  wire                pixelOut_ready;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_2_2_15;
  wire                pixelOut_payload_frame_line_endOfLine;
  wire                pixelOut_payload_frame_endOfFrame;
  wire                pixelOut_payload_endOfPack;
  reg                 pixel_videoOut_rValid;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_2_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_2_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_0_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_1_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_2_2_15;
  reg                 pixel_videoOut_rData_frame_line_endOfLine;
  reg                 pixel_videoOut_rData_frame_endOfFrame;
  reg                 pixel_videoOut_rData_endOfPack;
  wire                when_Stream_l342;
  wire                line_videoOut_m2sPipe_valid;
  wire                line_videoOut_m2sPipe_ready;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_0;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_1;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_2;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_3;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_4;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_5;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_6;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_7;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_8;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_9;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_10;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_11;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_12;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_13;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_14;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_15;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_0;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_1;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_2;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_3;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_4;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_5;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_6;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_7;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_8;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_9;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_10;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_11;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_12;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_13;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_14;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_15;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_0;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_1;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_2;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_3;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_4;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_5;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_6;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_7;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_8;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_9;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_10;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_11;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_12;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_13;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_14;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_2_15;
  wire                line_videoOut_m2sPipe_payload_frame_line_endOfLine;
  wire                line_videoOut_m2sPipe_payload_frame_endOfFrame;
  wire                line_videoOut_m2sPipe_payload_endOfPack;
  reg                 line_videoOut_rValid;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_0;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_1;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_2;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_3;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_4;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_5;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_6;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_7;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_8;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_9;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_10;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_11;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_12;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_13;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_14;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_15;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_0;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_1;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_2;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_3;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_4;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_5;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_6;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_7;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_8;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_9;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_10;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_11;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_12;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_13;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_14;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_15;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_0;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_1;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_2;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_3;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_4;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_5;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_6;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_7;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_8;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_9;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_10;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_11;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_12;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_13;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_14;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_2_15;
  reg                 line_videoOut_rData_frame_line_endOfLine;
  reg                 line_videoOut_rData_frame_endOfFrame;
  reg                 line_videoOut_rData_endOfPack;
  wire                when_Stream_l342_1;
  wire                line_videoOut_m2sPipe_s2mPipe_valid;
  wire                line_videoOut_m2sPipe_s2mPipe_ready;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_0;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_1;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_2;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_3;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_4;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_5;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_6;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_7;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_8;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_9;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_10;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_11;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_12;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_13;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_14;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_15;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_0;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_1;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_2;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_3;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_4;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_5;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_6;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_7;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_8;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_9;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_10;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_11;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_12;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_13;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_14;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_15;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_0;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_1;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_2;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_3;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_4;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_5;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_6;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_7;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_8;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_9;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_10;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_11;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_12;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_13;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_14;
  wire       [7:0]    line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_15;
  wire                line_videoOut_m2sPipe_s2mPipe_payload_frame_line_endOfLine;
  wire                line_videoOut_m2sPipe_s2mPipe_payload_frame_endOfFrame;
  wire                line_videoOut_m2sPipe_s2mPipe_payload_endOfPack;
  reg                 line_videoOut_m2sPipe_rValid;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_0;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_1;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_2;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_3;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_4;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_5;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_6;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_7;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_8;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_9;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_10;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_11;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_12;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_13;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_14;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_0_15;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_0;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_1;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_2;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_3;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_4;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_5;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_6;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_7;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_8;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_9;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_10;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_11;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_12;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_13;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_14;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_1_15;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_0;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_1;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_2;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_3;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_4;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_5;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_6;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_7;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_8;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_9;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_10;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_11;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_12;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_13;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_14;
  reg        [7:0]    line_videoOut_m2sPipe_rData_frame_line_pixel_2_15;
  reg                 line_videoOut_m2sPipe_rData_frame_line_endOfLine;
  reg                 line_videoOut_m2sPipe_rData_frame_endOfFrame;
  reg                 line_videoOut_m2sPipe_rData_endOfPack;

  LineBufferSame line (
    .videoIn_valid                             (videoIn_valid                                     ), //i
    .videoIn_ready                             (line_videoIn_ready                                ), //o
    .videoIn_payload_frame_line_pixel_0        (videoIn_payload_frame_line_pixel_0[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_1        (videoIn_payload_frame_line_pixel_1[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_2        (videoIn_payload_frame_line_pixel_2[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_3        (videoIn_payload_frame_line_pixel_3[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_4        (videoIn_payload_frame_line_pixel_4[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_5        (videoIn_payload_frame_line_pixel_5[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_6        (videoIn_payload_frame_line_pixel_6[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_7        (videoIn_payload_frame_line_pixel_7[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_8        (videoIn_payload_frame_line_pixel_8[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_9        (videoIn_payload_frame_line_pixel_9[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_10       (videoIn_payload_frame_line_pixel_10[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_11       (videoIn_payload_frame_line_pixel_11[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_12       (videoIn_payload_frame_line_pixel_12[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_13       (videoIn_payload_frame_line_pixel_13[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_14       (videoIn_payload_frame_line_pixel_14[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_15       (videoIn_payload_frame_line_pixel_15[7:0]          ), //i
    .videoIn_payload_frame_line_endOfLine      (videoIn_payload_frame_line_endOfLine              ), //i
    .videoIn_payload_frame_endOfFrame          (videoIn_payload_frame_endOfFrame                  ), //i
    .videoIn_payload_endOfPack                 (videoIn_payload_endOfPack                         ), //i
    .videoOut_valid                            (line_videoOut_valid                               ), //o
    .videoOut_ready                            (line_videoOut_ready                               ), //i
    .videoOut_payload_frame_line_pixel_0_0     (line_videoOut_payload_frame_line_pixel_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1     (line_videoOut_payload_frame_line_pixel_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2     (line_videoOut_payload_frame_line_pixel_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_3     (line_videoOut_payload_frame_line_pixel_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_4     (line_videoOut_payload_frame_line_pixel_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_5     (line_videoOut_payload_frame_line_pixel_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_6     (line_videoOut_payload_frame_line_pixel_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_7     (line_videoOut_payload_frame_line_pixel_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_8     (line_videoOut_payload_frame_line_pixel_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_9     (line_videoOut_payload_frame_line_pixel_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_10    (line_videoOut_payload_frame_line_pixel_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_11    (line_videoOut_payload_frame_line_pixel_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_12    (line_videoOut_payload_frame_line_pixel_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_13    (line_videoOut_payload_frame_line_pixel_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_14    (line_videoOut_payload_frame_line_pixel_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_15    (line_videoOut_payload_frame_line_pixel_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0     (line_videoOut_payload_frame_line_pixel_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1     (line_videoOut_payload_frame_line_pixel_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2     (line_videoOut_payload_frame_line_pixel_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_3     (line_videoOut_payload_frame_line_pixel_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_4     (line_videoOut_payload_frame_line_pixel_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_5     (line_videoOut_payload_frame_line_pixel_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_6     (line_videoOut_payload_frame_line_pixel_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_7     (line_videoOut_payload_frame_line_pixel_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_8     (line_videoOut_payload_frame_line_pixel_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_9     (line_videoOut_payload_frame_line_pixel_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_10    (line_videoOut_payload_frame_line_pixel_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_11    (line_videoOut_payload_frame_line_pixel_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_12    (line_videoOut_payload_frame_line_pixel_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_13    (line_videoOut_payload_frame_line_pixel_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_14    (line_videoOut_payload_frame_line_pixel_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_15    (line_videoOut_payload_frame_line_pixel_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_0     (line_videoOut_payload_frame_line_pixel_2_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_1     (line_videoOut_payload_frame_line_pixel_2_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_2     (line_videoOut_payload_frame_line_pixel_2_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_3     (line_videoOut_payload_frame_line_pixel_2_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_4     (line_videoOut_payload_frame_line_pixel_2_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_5     (line_videoOut_payload_frame_line_pixel_2_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_6     (line_videoOut_payload_frame_line_pixel_2_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_7     (line_videoOut_payload_frame_line_pixel_2_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_8     (line_videoOut_payload_frame_line_pixel_2_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_9     (line_videoOut_payload_frame_line_pixel_2_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_2_10    (line_videoOut_payload_frame_line_pixel_2_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_11    (line_videoOut_payload_frame_line_pixel_2_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_12    (line_videoOut_payload_frame_line_pixel_2_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_13    (line_videoOut_payload_frame_line_pixel_2_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_14    (line_videoOut_payload_frame_line_pixel_2_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_2_15    (line_videoOut_payload_frame_line_pixel_2_15[7:0]  ), //o
    .videoOut_payload_frame_line_endOfLine     (line_videoOut_payload_frame_line_endOfLine        ), //o
    .videoOut_payload_frame_endOfFrame         (line_videoOut_payload_frame_endOfFrame            ), //o
    .videoOut_payload_endOfPack                (line_videoOut_payload_endOfPack                   ), //o
    .clk                                       (clk                                               ), //i
    .reset                                     (reset                                             )  //i
  );
  PixelBufferSame pixel (
    .videoIn_valid                               (line_videoOut_m2sPipe_s2mPipe_valid                               ), //i
    .videoIn_ready                               (pixel_videoIn_ready                                               ), //o
    .videoIn_payload_frame_line_pixel_0_0        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_1        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_2        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_3        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_4        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_5        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_6        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_7        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_8        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_9        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_10       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_11       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_12       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_13       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_14       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_15       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_15[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_0        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_1        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_2        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_3        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_4        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_5        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_6        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_7        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_8        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_9        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_10       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_11       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_12       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_13       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_14       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_15       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_15[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_0        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_1        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_2        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_3        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_4        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_5        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_6        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_7        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_8        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_9        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_2_10       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_11       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_12       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_13       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_14       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_2_15       (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_15[7:0]  ), //i
    .videoIn_payload_frame_line_endOfLine        (line_videoOut_m2sPipe_s2mPipe_payload_frame_line_endOfLine        ), //i
    .videoIn_payload_frame_endOfFrame            (line_videoOut_m2sPipe_s2mPipe_payload_frame_endOfFrame            ), //i
    .videoIn_payload_endOfPack                   (line_videoOut_m2sPipe_s2mPipe_payload_endOfPack                   ), //i
    .videoOut_valid                              (pixel_videoOut_valid                                              ), //o
    .videoOut_ready                              (pixel_videoOut_ready                                              ), //i
    .videoOut_payload_frame_line_pixel_0_0_0     (pixel_videoOut_payload_frame_line_pixel_0_0_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_1     (pixel_videoOut_payload_frame_line_pixel_0_0_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_2     (pixel_videoOut_payload_frame_line_pixel_0_0_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_3     (pixel_videoOut_payload_frame_line_pixel_0_0_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_4     (pixel_videoOut_payload_frame_line_pixel_0_0_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_5     (pixel_videoOut_payload_frame_line_pixel_0_0_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_6     (pixel_videoOut_payload_frame_line_pixel_0_0_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_7     (pixel_videoOut_payload_frame_line_pixel_0_0_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_8     (pixel_videoOut_payload_frame_line_pixel_0_0_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_9     (pixel_videoOut_payload_frame_line_pixel_0_0_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_0_10    (pixel_videoOut_payload_frame_line_pixel_0_0_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_0_11    (pixel_videoOut_payload_frame_line_pixel_0_0_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_0_12    (pixel_videoOut_payload_frame_line_pixel_0_0_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_0_13    (pixel_videoOut_payload_frame_line_pixel_0_0_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_0_14    (pixel_videoOut_payload_frame_line_pixel_0_0_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_0_15    (pixel_videoOut_payload_frame_line_pixel_0_0_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_0     (pixel_videoOut_payload_frame_line_pixel_0_1_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_1     (pixel_videoOut_payload_frame_line_pixel_0_1_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_2     (pixel_videoOut_payload_frame_line_pixel_0_1_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_3     (pixel_videoOut_payload_frame_line_pixel_0_1_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_4     (pixel_videoOut_payload_frame_line_pixel_0_1_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_5     (pixel_videoOut_payload_frame_line_pixel_0_1_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_6     (pixel_videoOut_payload_frame_line_pixel_0_1_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_7     (pixel_videoOut_payload_frame_line_pixel_0_1_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_8     (pixel_videoOut_payload_frame_line_pixel_0_1_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_9     (pixel_videoOut_payload_frame_line_pixel_0_1_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_1_10    (pixel_videoOut_payload_frame_line_pixel_0_1_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_11    (pixel_videoOut_payload_frame_line_pixel_0_1_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_12    (pixel_videoOut_payload_frame_line_pixel_0_1_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_13    (pixel_videoOut_payload_frame_line_pixel_0_1_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_14    (pixel_videoOut_payload_frame_line_pixel_0_1_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_1_15    (pixel_videoOut_payload_frame_line_pixel_0_1_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_0     (pixel_videoOut_payload_frame_line_pixel_0_2_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_1     (pixel_videoOut_payload_frame_line_pixel_0_2_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_2     (pixel_videoOut_payload_frame_line_pixel_0_2_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_3     (pixel_videoOut_payload_frame_line_pixel_0_2_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_4     (pixel_videoOut_payload_frame_line_pixel_0_2_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_5     (pixel_videoOut_payload_frame_line_pixel_0_2_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_6     (pixel_videoOut_payload_frame_line_pixel_0_2_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_7     (pixel_videoOut_payload_frame_line_pixel_0_2_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_8     (pixel_videoOut_payload_frame_line_pixel_0_2_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_9     (pixel_videoOut_payload_frame_line_pixel_0_2_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_0_2_10    (pixel_videoOut_payload_frame_line_pixel_0_2_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_11    (pixel_videoOut_payload_frame_line_pixel_0_2_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_12    (pixel_videoOut_payload_frame_line_pixel_0_2_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_13    (pixel_videoOut_payload_frame_line_pixel_0_2_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_14    (pixel_videoOut_payload_frame_line_pixel_0_2_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_0_2_15    (pixel_videoOut_payload_frame_line_pixel_0_2_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_0     (pixel_videoOut_payload_frame_line_pixel_1_0_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_1     (pixel_videoOut_payload_frame_line_pixel_1_0_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_2     (pixel_videoOut_payload_frame_line_pixel_1_0_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_3     (pixel_videoOut_payload_frame_line_pixel_1_0_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_4     (pixel_videoOut_payload_frame_line_pixel_1_0_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_5     (pixel_videoOut_payload_frame_line_pixel_1_0_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_6     (pixel_videoOut_payload_frame_line_pixel_1_0_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_7     (pixel_videoOut_payload_frame_line_pixel_1_0_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_8     (pixel_videoOut_payload_frame_line_pixel_1_0_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_9     (pixel_videoOut_payload_frame_line_pixel_1_0_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_0_10    (pixel_videoOut_payload_frame_line_pixel_1_0_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_11    (pixel_videoOut_payload_frame_line_pixel_1_0_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_12    (pixel_videoOut_payload_frame_line_pixel_1_0_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_13    (pixel_videoOut_payload_frame_line_pixel_1_0_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_14    (pixel_videoOut_payload_frame_line_pixel_1_0_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_0_15    (pixel_videoOut_payload_frame_line_pixel_1_0_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_0     (pixel_videoOut_payload_frame_line_pixel_1_1_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_1     (pixel_videoOut_payload_frame_line_pixel_1_1_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_2     (pixel_videoOut_payload_frame_line_pixel_1_1_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_3     (pixel_videoOut_payload_frame_line_pixel_1_1_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_4     (pixel_videoOut_payload_frame_line_pixel_1_1_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_5     (pixel_videoOut_payload_frame_line_pixel_1_1_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_6     (pixel_videoOut_payload_frame_line_pixel_1_1_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_7     (pixel_videoOut_payload_frame_line_pixel_1_1_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_8     (pixel_videoOut_payload_frame_line_pixel_1_1_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_9     (pixel_videoOut_payload_frame_line_pixel_1_1_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_1_10    (pixel_videoOut_payload_frame_line_pixel_1_1_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_11    (pixel_videoOut_payload_frame_line_pixel_1_1_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_12    (pixel_videoOut_payload_frame_line_pixel_1_1_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_13    (pixel_videoOut_payload_frame_line_pixel_1_1_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_14    (pixel_videoOut_payload_frame_line_pixel_1_1_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_1_15    (pixel_videoOut_payload_frame_line_pixel_1_1_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_0     (pixel_videoOut_payload_frame_line_pixel_1_2_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_1     (pixel_videoOut_payload_frame_line_pixel_1_2_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_2     (pixel_videoOut_payload_frame_line_pixel_1_2_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_3     (pixel_videoOut_payload_frame_line_pixel_1_2_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_4     (pixel_videoOut_payload_frame_line_pixel_1_2_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_5     (pixel_videoOut_payload_frame_line_pixel_1_2_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_6     (pixel_videoOut_payload_frame_line_pixel_1_2_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_7     (pixel_videoOut_payload_frame_line_pixel_1_2_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_8     (pixel_videoOut_payload_frame_line_pixel_1_2_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_9     (pixel_videoOut_payload_frame_line_pixel_1_2_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_1_2_10    (pixel_videoOut_payload_frame_line_pixel_1_2_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_11    (pixel_videoOut_payload_frame_line_pixel_1_2_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_12    (pixel_videoOut_payload_frame_line_pixel_1_2_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_13    (pixel_videoOut_payload_frame_line_pixel_1_2_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_14    (pixel_videoOut_payload_frame_line_pixel_1_2_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_1_2_15    (pixel_videoOut_payload_frame_line_pixel_1_2_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_0     (pixel_videoOut_payload_frame_line_pixel_2_0_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_1     (pixel_videoOut_payload_frame_line_pixel_2_0_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_2     (pixel_videoOut_payload_frame_line_pixel_2_0_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_3     (pixel_videoOut_payload_frame_line_pixel_2_0_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_4     (pixel_videoOut_payload_frame_line_pixel_2_0_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_5     (pixel_videoOut_payload_frame_line_pixel_2_0_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_6     (pixel_videoOut_payload_frame_line_pixel_2_0_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_7     (pixel_videoOut_payload_frame_line_pixel_2_0_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_8     (pixel_videoOut_payload_frame_line_pixel_2_0_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_9     (pixel_videoOut_payload_frame_line_pixel_2_0_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_0_10    (pixel_videoOut_payload_frame_line_pixel_2_0_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_11    (pixel_videoOut_payload_frame_line_pixel_2_0_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_12    (pixel_videoOut_payload_frame_line_pixel_2_0_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_13    (pixel_videoOut_payload_frame_line_pixel_2_0_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_14    (pixel_videoOut_payload_frame_line_pixel_2_0_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_0_15    (pixel_videoOut_payload_frame_line_pixel_2_0_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_0     (pixel_videoOut_payload_frame_line_pixel_2_1_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_1     (pixel_videoOut_payload_frame_line_pixel_2_1_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_2     (pixel_videoOut_payload_frame_line_pixel_2_1_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_3     (pixel_videoOut_payload_frame_line_pixel_2_1_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_4     (pixel_videoOut_payload_frame_line_pixel_2_1_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_5     (pixel_videoOut_payload_frame_line_pixel_2_1_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_6     (pixel_videoOut_payload_frame_line_pixel_2_1_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_7     (pixel_videoOut_payload_frame_line_pixel_2_1_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_8     (pixel_videoOut_payload_frame_line_pixel_2_1_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_9     (pixel_videoOut_payload_frame_line_pixel_2_1_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_1_10    (pixel_videoOut_payload_frame_line_pixel_2_1_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_11    (pixel_videoOut_payload_frame_line_pixel_2_1_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_12    (pixel_videoOut_payload_frame_line_pixel_2_1_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_13    (pixel_videoOut_payload_frame_line_pixel_2_1_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_14    (pixel_videoOut_payload_frame_line_pixel_2_1_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_1_15    (pixel_videoOut_payload_frame_line_pixel_2_1_15[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_0     (pixel_videoOut_payload_frame_line_pixel_2_2_0[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_1     (pixel_videoOut_payload_frame_line_pixel_2_2_1[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_2     (pixel_videoOut_payload_frame_line_pixel_2_2_2[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_3     (pixel_videoOut_payload_frame_line_pixel_2_2_3[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_4     (pixel_videoOut_payload_frame_line_pixel_2_2_4[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_5     (pixel_videoOut_payload_frame_line_pixel_2_2_5[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_6     (pixel_videoOut_payload_frame_line_pixel_2_2_6[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_7     (pixel_videoOut_payload_frame_line_pixel_2_2_7[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_8     (pixel_videoOut_payload_frame_line_pixel_2_2_8[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_9     (pixel_videoOut_payload_frame_line_pixel_2_2_9[7:0]                ), //o
    .videoOut_payload_frame_line_pixel_2_2_10    (pixel_videoOut_payload_frame_line_pixel_2_2_10[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_11    (pixel_videoOut_payload_frame_line_pixel_2_2_11[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_12    (pixel_videoOut_payload_frame_line_pixel_2_2_12[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_13    (pixel_videoOut_payload_frame_line_pixel_2_2_13[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_14    (pixel_videoOut_payload_frame_line_pixel_2_2_14[7:0]               ), //o
    .videoOut_payload_frame_line_pixel_2_2_15    (pixel_videoOut_payload_frame_line_pixel_2_2_15[7:0]               ), //o
    .videoOut_payload_frame_line_endOfLine       (pixel_videoOut_payload_frame_line_endOfLine                       ), //o
    .videoOut_payload_frame_endOfFrame           (pixel_videoOut_payload_frame_endOfFrame                           ), //o
    .videoOut_payload_endOfPack                  (pixel_videoOut_payload_endOfPack                                  ), //o
    .clk                                         (clk                                                               ), //i
    .reset                                       (reset                                                             )  //i
  );
  always @(*) begin
    pixel_videoOut_ready = pixelOut_ready;
    if(when_Stream_l342) begin
      pixel_videoOut_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! pixelOut_valid);
  assign pixelOut_valid = pixel_videoOut_rValid;
  assign pixelOut_payload_frame_line_pixel_0_0_0 = pixel_videoOut_rData_frame_line_pixel_0_0_0;
  assign pixelOut_payload_frame_line_pixel_0_0_1 = pixel_videoOut_rData_frame_line_pixel_0_0_1;
  assign pixelOut_payload_frame_line_pixel_0_0_2 = pixel_videoOut_rData_frame_line_pixel_0_0_2;
  assign pixelOut_payload_frame_line_pixel_0_0_3 = pixel_videoOut_rData_frame_line_pixel_0_0_3;
  assign pixelOut_payload_frame_line_pixel_0_0_4 = pixel_videoOut_rData_frame_line_pixel_0_0_4;
  assign pixelOut_payload_frame_line_pixel_0_0_5 = pixel_videoOut_rData_frame_line_pixel_0_0_5;
  assign pixelOut_payload_frame_line_pixel_0_0_6 = pixel_videoOut_rData_frame_line_pixel_0_0_6;
  assign pixelOut_payload_frame_line_pixel_0_0_7 = pixel_videoOut_rData_frame_line_pixel_0_0_7;
  assign pixelOut_payload_frame_line_pixel_0_0_8 = pixel_videoOut_rData_frame_line_pixel_0_0_8;
  assign pixelOut_payload_frame_line_pixel_0_0_9 = pixel_videoOut_rData_frame_line_pixel_0_0_9;
  assign pixelOut_payload_frame_line_pixel_0_0_10 = pixel_videoOut_rData_frame_line_pixel_0_0_10;
  assign pixelOut_payload_frame_line_pixel_0_0_11 = pixel_videoOut_rData_frame_line_pixel_0_0_11;
  assign pixelOut_payload_frame_line_pixel_0_0_12 = pixel_videoOut_rData_frame_line_pixel_0_0_12;
  assign pixelOut_payload_frame_line_pixel_0_0_13 = pixel_videoOut_rData_frame_line_pixel_0_0_13;
  assign pixelOut_payload_frame_line_pixel_0_0_14 = pixel_videoOut_rData_frame_line_pixel_0_0_14;
  assign pixelOut_payload_frame_line_pixel_0_0_15 = pixel_videoOut_rData_frame_line_pixel_0_0_15;
  assign pixelOut_payload_frame_line_pixel_0_1_0 = pixel_videoOut_rData_frame_line_pixel_0_1_0;
  assign pixelOut_payload_frame_line_pixel_0_1_1 = pixel_videoOut_rData_frame_line_pixel_0_1_1;
  assign pixelOut_payload_frame_line_pixel_0_1_2 = pixel_videoOut_rData_frame_line_pixel_0_1_2;
  assign pixelOut_payload_frame_line_pixel_0_1_3 = pixel_videoOut_rData_frame_line_pixel_0_1_3;
  assign pixelOut_payload_frame_line_pixel_0_1_4 = pixel_videoOut_rData_frame_line_pixel_0_1_4;
  assign pixelOut_payload_frame_line_pixel_0_1_5 = pixel_videoOut_rData_frame_line_pixel_0_1_5;
  assign pixelOut_payload_frame_line_pixel_0_1_6 = pixel_videoOut_rData_frame_line_pixel_0_1_6;
  assign pixelOut_payload_frame_line_pixel_0_1_7 = pixel_videoOut_rData_frame_line_pixel_0_1_7;
  assign pixelOut_payload_frame_line_pixel_0_1_8 = pixel_videoOut_rData_frame_line_pixel_0_1_8;
  assign pixelOut_payload_frame_line_pixel_0_1_9 = pixel_videoOut_rData_frame_line_pixel_0_1_9;
  assign pixelOut_payload_frame_line_pixel_0_1_10 = pixel_videoOut_rData_frame_line_pixel_0_1_10;
  assign pixelOut_payload_frame_line_pixel_0_1_11 = pixel_videoOut_rData_frame_line_pixel_0_1_11;
  assign pixelOut_payload_frame_line_pixel_0_1_12 = pixel_videoOut_rData_frame_line_pixel_0_1_12;
  assign pixelOut_payload_frame_line_pixel_0_1_13 = pixel_videoOut_rData_frame_line_pixel_0_1_13;
  assign pixelOut_payload_frame_line_pixel_0_1_14 = pixel_videoOut_rData_frame_line_pixel_0_1_14;
  assign pixelOut_payload_frame_line_pixel_0_1_15 = pixel_videoOut_rData_frame_line_pixel_0_1_15;
  assign pixelOut_payload_frame_line_pixel_0_2_0 = pixel_videoOut_rData_frame_line_pixel_0_2_0;
  assign pixelOut_payload_frame_line_pixel_0_2_1 = pixel_videoOut_rData_frame_line_pixel_0_2_1;
  assign pixelOut_payload_frame_line_pixel_0_2_2 = pixel_videoOut_rData_frame_line_pixel_0_2_2;
  assign pixelOut_payload_frame_line_pixel_0_2_3 = pixel_videoOut_rData_frame_line_pixel_0_2_3;
  assign pixelOut_payload_frame_line_pixel_0_2_4 = pixel_videoOut_rData_frame_line_pixel_0_2_4;
  assign pixelOut_payload_frame_line_pixel_0_2_5 = pixel_videoOut_rData_frame_line_pixel_0_2_5;
  assign pixelOut_payload_frame_line_pixel_0_2_6 = pixel_videoOut_rData_frame_line_pixel_0_2_6;
  assign pixelOut_payload_frame_line_pixel_0_2_7 = pixel_videoOut_rData_frame_line_pixel_0_2_7;
  assign pixelOut_payload_frame_line_pixel_0_2_8 = pixel_videoOut_rData_frame_line_pixel_0_2_8;
  assign pixelOut_payload_frame_line_pixel_0_2_9 = pixel_videoOut_rData_frame_line_pixel_0_2_9;
  assign pixelOut_payload_frame_line_pixel_0_2_10 = pixel_videoOut_rData_frame_line_pixel_0_2_10;
  assign pixelOut_payload_frame_line_pixel_0_2_11 = pixel_videoOut_rData_frame_line_pixel_0_2_11;
  assign pixelOut_payload_frame_line_pixel_0_2_12 = pixel_videoOut_rData_frame_line_pixel_0_2_12;
  assign pixelOut_payload_frame_line_pixel_0_2_13 = pixel_videoOut_rData_frame_line_pixel_0_2_13;
  assign pixelOut_payload_frame_line_pixel_0_2_14 = pixel_videoOut_rData_frame_line_pixel_0_2_14;
  assign pixelOut_payload_frame_line_pixel_0_2_15 = pixel_videoOut_rData_frame_line_pixel_0_2_15;
  assign pixelOut_payload_frame_line_pixel_1_0_0 = pixel_videoOut_rData_frame_line_pixel_1_0_0;
  assign pixelOut_payload_frame_line_pixel_1_0_1 = pixel_videoOut_rData_frame_line_pixel_1_0_1;
  assign pixelOut_payload_frame_line_pixel_1_0_2 = pixel_videoOut_rData_frame_line_pixel_1_0_2;
  assign pixelOut_payload_frame_line_pixel_1_0_3 = pixel_videoOut_rData_frame_line_pixel_1_0_3;
  assign pixelOut_payload_frame_line_pixel_1_0_4 = pixel_videoOut_rData_frame_line_pixel_1_0_4;
  assign pixelOut_payload_frame_line_pixel_1_0_5 = pixel_videoOut_rData_frame_line_pixel_1_0_5;
  assign pixelOut_payload_frame_line_pixel_1_0_6 = pixel_videoOut_rData_frame_line_pixel_1_0_6;
  assign pixelOut_payload_frame_line_pixel_1_0_7 = pixel_videoOut_rData_frame_line_pixel_1_0_7;
  assign pixelOut_payload_frame_line_pixel_1_0_8 = pixel_videoOut_rData_frame_line_pixel_1_0_8;
  assign pixelOut_payload_frame_line_pixel_1_0_9 = pixel_videoOut_rData_frame_line_pixel_1_0_9;
  assign pixelOut_payload_frame_line_pixel_1_0_10 = pixel_videoOut_rData_frame_line_pixel_1_0_10;
  assign pixelOut_payload_frame_line_pixel_1_0_11 = pixel_videoOut_rData_frame_line_pixel_1_0_11;
  assign pixelOut_payload_frame_line_pixel_1_0_12 = pixel_videoOut_rData_frame_line_pixel_1_0_12;
  assign pixelOut_payload_frame_line_pixel_1_0_13 = pixel_videoOut_rData_frame_line_pixel_1_0_13;
  assign pixelOut_payload_frame_line_pixel_1_0_14 = pixel_videoOut_rData_frame_line_pixel_1_0_14;
  assign pixelOut_payload_frame_line_pixel_1_0_15 = pixel_videoOut_rData_frame_line_pixel_1_0_15;
  assign pixelOut_payload_frame_line_pixel_1_1_0 = pixel_videoOut_rData_frame_line_pixel_1_1_0;
  assign pixelOut_payload_frame_line_pixel_1_1_1 = pixel_videoOut_rData_frame_line_pixel_1_1_1;
  assign pixelOut_payload_frame_line_pixel_1_1_2 = pixel_videoOut_rData_frame_line_pixel_1_1_2;
  assign pixelOut_payload_frame_line_pixel_1_1_3 = pixel_videoOut_rData_frame_line_pixel_1_1_3;
  assign pixelOut_payload_frame_line_pixel_1_1_4 = pixel_videoOut_rData_frame_line_pixel_1_1_4;
  assign pixelOut_payload_frame_line_pixel_1_1_5 = pixel_videoOut_rData_frame_line_pixel_1_1_5;
  assign pixelOut_payload_frame_line_pixel_1_1_6 = pixel_videoOut_rData_frame_line_pixel_1_1_6;
  assign pixelOut_payload_frame_line_pixel_1_1_7 = pixel_videoOut_rData_frame_line_pixel_1_1_7;
  assign pixelOut_payload_frame_line_pixel_1_1_8 = pixel_videoOut_rData_frame_line_pixel_1_1_8;
  assign pixelOut_payload_frame_line_pixel_1_1_9 = pixel_videoOut_rData_frame_line_pixel_1_1_9;
  assign pixelOut_payload_frame_line_pixel_1_1_10 = pixel_videoOut_rData_frame_line_pixel_1_1_10;
  assign pixelOut_payload_frame_line_pixel_1_1_11 = pixel_videoOut_rData_frame_line_pixel_1_1_11;
  assign pixelOut_payload_frame_line_pixel_1_1_12 = pixel_videoOut_rData_frame_line_pixel_1_1_12;
  assign pixelOut_payload_frame_line_pixel_1_1_13 = pixel_videoOut_rData_frame_line_pixel_1_1_13;
  assign pixelOut_payload_frame_line_pixel_1_1_14 = pixel_videoOut_rData_frame_line_pixel_1_1_14;
  assign pixelOut_payload_frame_line_pixel_1_1_15 = pixel_videoOut_rData_frame_line_pixel_1_1_15;
  assign pixelOut_payload_frame_line_pixel_1_2_0 = pixel_videoOut_rData_frame_line_pixel_1_2_0;
  assign pixelOut_payload_frame_line_pixel_1_2_1 = pixel_videoOut_rData_frame_line_pixel_1_2_1;
  assign pixelOut_payload_frame_line_pixel_1_2_2 = pixel_videoOut_rData_frame_line_pixel_1_2_2;
  assign pixelOut_payload_frame_line_pixel_1_2_3 = pixel_videoOut_rData_frame_line_pixel_1_2_3;
  assign pixelOut_payload_frame_line_pixel_1_2_4 = pixel_videoOut_rData_frame_line_pixel_1_2_4;
  assign pixelOut_payload_frame_line_pixel_1_2_5 = pixel_videoOut_rData_frame_line_pixel_1_2_5;
  assign pixelOut_payload_frame_line_pixel_1_2_6 = pixel_videoOut_rData_frame_line_pixel_1_2_6;
  assign pixelOut_payload_frame_line_pixel_1_2_7 = pixel_videoOut_rData_frame_line_pixel_1_2_7;
  assign pixelOut_payload_frame_line_pixel_1_2_8 = pixel_videoOut_rData_frame_line_pixel_1_2_8;
  assign pixelOut_payload_frame_line_pixel_1_2_9 = pixel_videoOut_rData_frame_line_pixel_1_2_9;
  assign pixelOut_payload_frame_line_pixel_1_2_10 = pixel_videoOut_rData_frame_line_pixel_1_2_10;
  assign pixelOut_payload_frame_line_pixel_1_2_11 = pixel_videoOut_rData_frame_line_pixel_1_2_11;
  assign pixelOut_payload_frame_line_pixel_1_2_12 = pixel_videoOut_rData_frame_line_pixel_1_2_12;
  assign pixelOut_payload_frame_line_pixel_1_2_13 = pixel_videoOut_rData_frame_line_pixel_1_2_13;
  assign pixelOut_payload_frame_line_pixel_1_2_14 = pixel_videoOut_rData_frame_line_pixel_1_2_14;
  assign pixelOut_payload_frame_line_pixel_1_2_15 = pixel_videoOut_rData_frame_line_pixel_1_2_15;
  assign pixelOut_payload_frame_line_pixel_2_0_0 = pixel_videoOut_rData_frame_line_pixel_2_0_0;
  assign pixelOut_payload_frame_line_pixel_2_0_1 = pixel_videoOut_rData_frame_line_pixel_2_0_1;
  assign pixelOut_payload_frame_line_pixel_2_0_2 = pixel_videoOut_rData_frame_line_pixel_2_0_2;
  assign pixelOut_payload_frame_line_pixel_2_0_3 = pixel_videoOut_rData_frame_line_pixel_2_0_3;
  assign pixelOut_payload_frame_line_pixel_2_0_4 = pixel_videoOut_rData_frame_line_pixel_2_0_4;
  assign pixelOut_payload_frame_line_pixel_2_0_5 = pixel_videoOut_rData_frame_line_pixel_2_0_5;
  assign pixelOut_payload_frame_line_pixel_2_0_6 = pixel_videoOut_rData_frame_line_pixel_2_0_6;
  assign pixelOut_payload_frame_line_pixel_2_0_7 = pixel_videoOut_rData_frame_line_pixel_2_0_7;
  assign pixelOut_payload_frame_line_pixel_2_0_8 = pixel_videoOut_rData_frame_line_pixel_2_0_8;
  assign pixelOut_payload_frame_line_pixel_2_0_9 = pixel_videoOut_rData_frame_line_pixel_2_0_9;
  assign pixelOut_payload_frame_line_pixel_2_0_10 = pixel_videoOut_rData_frame_line_pixel_2_0_10;
  assign pixelOut_payload_frame_line_pixel_2_0_11 = pixel_videoOut_rData_frame_line_pixel_2_0_11;
  assign pixelOut_payload_frame_line_pixel_2_0_12 = pixel_videoOut_rData_frame_line_pixel_2_0_12;
  assign pixelOut_payload_frame_line_pixel_2_0_13 = pixel_videoOut_rData_frame_line_pixel_2_0_13;
  assign pixelOut_payload_frame_line_pixel_2_0_14 = pixel_videoOut_rData_frame_line_pixel_2_0_14;
  assign pixelOut_payload_frame_line_pixel_2_0_15 = pixel_videoOut_rData_frame_line_pixel_2_0_15;
  assign pixelOut_payload_frame_line_pixel_2_1_0 = pixel_videoOut_rData_frame_line_pixel_2_1_0;
  assign pixelOut_payload_frame_line_pixel_2_1_1 = pixel_videoOut_rData_frame_line_pixel_2_1_1;
  assign pixelOut_payload_frame_line_pixel_2_1_2 = pixel_videoOut_rData_frame_line_pixel_2_1_2;
  assign pixelOut_payload_frame_line_pixel_2_1_3 = pixel_videoOut_rData_frame_line_pixel_2_1_3;
  assign pixelOut_payload_frame_line_pixel_2_1_4 = pixel_videoOut_rData_frame_line_pixel_2_1_4;
  assign pixelOut_payload_frame_line_pixel_2_1_5 = pixel_videoOut_rData_frame_line_pixel_2_1_5;
  assign pixelOut_payload_frame_line_pixel_2_1_6 = pixel_videoOut_rData_frame_line_pixel_2_1_6;
  assign pixelOut_payload_frame_line_pixel_2_1_7 = pixel_videoOut_rData_frame_line_pixel_2_1_7;
  assign pixelOut_payload_frame_line_pixel_2_1_8 = pixel_videoOut_rData_frame_line_pixel_2_1_8;
  assign pixelOut_payload_frame_line_pixel_2_1_9 = pixel_videoOut_rData_frame_line_pixel_2_1_9;
  assign pixelOut_payload_frame_line_pixel_2_1_10 = pixel_videoOut_rData_frame_line_pixel_2_1_10;
  assign pixelOut_payload_frame_line_pixel_2_1_11 = pixel_videoOut_rData_frame_line_pixel_2_1_11;
  assign pixelOut_payload_frame_line_pixel_2_1_12 = pixel_videoOut_rData_frame_line_pixel_2_1_12;
  assign pixelOut_payload_frame_line_pixel_2_1_13 = pixel_videoOut_rData_frame_line_pixel_2_1_13;
  assign pixelOut_payload_frame_line_pixel_2_1_14 = pixel_videoOut_rData_frame_line_pixel_2_1_14;
  assign pixelOut_payload_frame_line_pixel_2_1_15 = pixel_videoOut_rData_frame_line_pixel_2_1_15;
  assign pixelOut_payload_frame_line_pixel_2_2_0 = pixel_videoOut_rData_frame_line_pixel_2_2_0;
  assign pixelOut_payload_frame_line_pixel_2_2_1 = pixel_videoOut_rData_frame_line_pixel_2_2_1;
  assign pixelOut_payload_frame_line_pixel_2_2_2 = pixel_videoOut_rData_frame_line_pixel_2_2_2;
  assign pixelOut_payload_frame_line_pixel_2_2_3 = pixel_videoOut_rData_frame_line_pixel_2_2_3;
  assign pixelOut_payload_frame_line_pixel_2_2_4 = pixel_videoOut_rData_frame_line_pixel_2_2_4;
  assign pixelOut_payload_frame_line_pixel_2_2_5 = pixel_videoOut_rData_frame_line_pixel_2_2_5;
  assign pixelOut_payload_frame_line_pixel_2_2_6 = pixel_videoOut_rData_frame_line_pixel_2_2_6;
  assign pixelOut_payload_frame_line_pixel_2_2_7 = pixel_videoOut_rData_frame_line_pixel_2_2_7;
  assign pixelOut_payload_frame_line_pixel_2_2_8 = pixel_videoOut_rData_frame_line_pixel_2_2_8;
  assign pixelOut_payload_frame_line_pixel_2_2_9 = pixel_videoOut_rData_frame_line_pixel_2_2_9;
  assign pixelOut_payload_frame_line_pixel_2_2_10 = pixel_videoOut_rData_frame_line_pixel_2_2_10;
  assign pixelOut_payload_frame_line_pixel_2_2_11 = pixel_videoOut_rData_frame_line_pixel_2_2_11;
  assign pixelOut_payload_frame_line_pixel_2_2_12 = pixel_videoOut_rData_frame_line_pixel_2_2_12;
  assign pixelOut_payload_frame_line_pixel_2_2_13 = pixel_videoOut_rData_frame_line_pixel_2_2_13;
  assign pixelOut_payload_frame_line_pixel_2_2_14 = pixel_videoOut_rData_frame_line_pixel_2_2_14;
  assign pixelOut_payload_frame_line_pixel_2_2_15 = pixel_videoOut_rData_frame_line_pixel_2_2_15;
  assign pixelOut_payload_frame_line_endOfLine = pixel_videoOut_rData_frame_line_endOfLine;
  assign pixelOut_payload_frame_endOfFrame = pixel_videoOut_rData_frame_endOfFrame;
  assign pixelOut_payload_endOfPack = pixel_videoOut_rData_endOfPack;
  assign videoIn_ready = line_videoIn_ready;
  always @(*) begin
    line_videoOut_ready = line_videoOut_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      line_videoOut_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! line_videoOut_m2sPipe_valid);
  assign line_videoOut_m2sPipe_valid = line_videoOut_rValid;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_0 = line_videoOut_rData_frame_line_pixel_0_0;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_1 = line_videoOut_rData_frame_line_pixel_0_1;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_2 = line_videoOut_rData_frame_line_pixel_0_2;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_3 = line_videoOut_rData_frame_line_pixel_0_3;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_4 = line_videoOut_rData_frame_line_pixel_0_4;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_5 = line_videoOut_rData_frame_line_pixel_0_5;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_6 = line_videoOut_rData_frame_line_pixel_0_6;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_7 = line_videoOut_rData_frame_line_pixel_0_7;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_8 = line_videoOut_rData_frame_line_pixel_0_8;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_9 = line_videoOut_rData_frame_line_pixel_0_9;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_10 = line_videoOut_rData_frame_line_pixel_0_10;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_11 = line_videoOut_rData_frame_line_pixel_0_11;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_12 = line_videoOut_rData_frame_line_pixel_0_12;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_13 = line_videoOut_rData_frame_line_pixel_0_13;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_14 = line_videoOut_rData_frame_line_pixel_0_14;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_15 = line_videoOut_rData_frame_line_pixel_0_15;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_0 = line_videoOut_rData_frame_line_pixel_1_0;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_1 = line_videoOut_rData_frame_line_pixel_1_1;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_2 = line_videoOut_rData_frame_line_pixel_1_2;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_3 = line_videoOut_rData_frame_line_pixel_1_3;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_4 = line_videoOut_rData_frame_line_pixel_1_4;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_5 = line_videoOut_rData_frame_line_pixel_1_5;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_6 = line_videoOut_rData_frame_line_pixel_1_6;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_7 = line_videoOut_rData_frame_line_pixel_1_7;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_8 = line_videoOut_rData_frame_line_pixel_1_8;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_9 = line_videoOut_rData_frame_line_pixel_1_9;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_10 = line_videoOut_rData_frame_line_pixel_1_10;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_11 = line_videoOut_rData_frame_line_pixel_1_11;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_12 = line_videoOut_rData_frame_line_pixel_1_12;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_13 = line_videoOut_rData_frame_line_pixel_1_13;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_14 = line_videoOut_rData_frame_line_pixel_1_14;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_15 = line_videoOut_rData_frame_line_pixel_1_15;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_0 = line_videoOut_rData_frame_line_pixel_2_0;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_1 = line_videoOut_rData_frame_line_pixel_2_1;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_2 = line_videoOut_rData_frame_line_pixel_2_2;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_3 = line_videoOut_rData_frame_line_pixel_2_3;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_4 = line_videoOut_rData_frame_line_pixel_2_4;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_5 = line_videoOut_rData_frame_line_pixel_2_5;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_6 = line_videoOut_rData_frame_line_pixel_2_6;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_7 = line_videoOut_rData_frame_line_pixel_2_7;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_8 = line_videoOut_rData_frame_line_pixel_2_8;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_9 = line_videoOut_rData_frame_line_pixel_2_9;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_10 = line_videoOut_rData_frame_line_pixel_2_10;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_11 = line_videoOut_rData_frame_line_pixel_2_11;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_12 = line_videoOut_rData_frame_line_pixel_2_12;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_13 = line_videoOut_rData_frame_line_pixel_2_13;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_14 = line_videoOut_rData_frame_line_pixel_2_14;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_2_15 = line_videoOut_rData_frame_line_pixel_2_15;
  assign line_videoOut_m2sPipe_payload_frame_line_endOfLine = line_videoOut_rData_frame_line_endOfLine;
  assign line_videoOut_m2sPipe_payload_frame_endOfFrame = line_videoOut_rData_frame_endOfFrame;
  assign line_videoOut_m2sPipe_payload_endOfPack = line_videoOut_rData_endOfPack;
  assign line_videoOut_m2sPipe_ready = (! line_videoOut_m2sPipe_rValid);
  assign line_videoOut_m2sPipe_s2mPipe_valid = (line_videoOut_m2sPipe_valid || line_videoOut_m2sPipe_rValid);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_0 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_0 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_0);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_1 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_1 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_1);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_2 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_2 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_2);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_3 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_3 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_3);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_4 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_4 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_4);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_5 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_5 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_5);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_6 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_6 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_6);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_7 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_7 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_7);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_8 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_8 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_8);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_9 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_9 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_9);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_10 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_10 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_10);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_11 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_11 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_11);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_12 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_12 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_12);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_13 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_13 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_13);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_14 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_14 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_14);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_0_15 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_0_15 : line_videoOut_m2sPipe_payload_frame_line_pixel_0_15);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_0 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_0 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_0);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_1 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_1 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_1);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_2 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_2 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_2);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_3 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_3 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_3);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_4 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_4 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_4);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_5 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_5 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_5);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_6 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_6 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_6);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_7 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_7 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_7);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_8 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_8 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_8);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_9 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_9 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_9);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_10 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_10 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_10);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_11 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_11 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_11);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_12 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_12 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_12);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_13 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_13 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_13);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_14 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_14 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_14);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_1_15 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_1_15 : line_videoOut_m2sPipe_payload_frame_line_pixel_1_15);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_0 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_0 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_0);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_1 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_1 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_1);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_2 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_2 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_2);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_3 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_3 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_3);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_4 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_4 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_4);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_5 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_5 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_5);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_6 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_6 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_6);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_7 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_7 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_7);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_8 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_8 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_8);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_9 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_9 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_9);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_10 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_10 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_10);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_11 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_11 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_11);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_12 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_12 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_12);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_13 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_13 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_13);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_14 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_14 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_14);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_pixel_2_15 = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_pixel_2_15 : line_videoOut_m2sPipe_payload_frame_line_pixel_2_15);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_line_endOfLine = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_line_endOfLine : line_videoOut_m2sPipe_payload_frame_line_endOfLine);
  assign line_videoOut_m2sPipe_s2mPipe_payload_frame_endOfFrame = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_frame_endOfFrame : line_videoOut_m2sPipe_payload_frame_endOfFrame);
  assign line_videoOut_m2sPipe_s2mPipe_payload_endOfPack = (line_videoOut_m2sPipe_rValid ? line_videoOut_m2sPipe_rData_endOfPack : line_videoOut_m2sPipe_payload_endOfPack);
  assign line_videoOut_m2sPipe_s2mPipe_ready = pixel_videoIn_ready;
  assign videoOut_valid = pixelOut_valid;
  assign pixelOut_ready = videoOut_ready;
  assign videoOut_payload_endOfPack = pixelOut_payload_endOfPack;
  assign videoOut_payload_frame_endOfFrame = pixelOut_payload_frame_endOfFrame;
  assign videoOut_payload_frame_line_endOfLine = pixelOut_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_line_pixel_0_0_0 = pixelOut_payload_frame_line_pixel_0_0_0;
  assign videoOut_payload_frame_line_pixel_0_0_1 = pixelOut_payload_frame_line_pixel_0_0_1;
  assign videoOut_payload_frame_line_pixel_0_0_2 = pixelOut_payload_frame_line_pixel_0_0_2;
  assign videoOut_payload_frame_line_pixel_0_0_3 = pixelOut_payload_frame_line_pixel_0_0_3;
  assign videoOut_payload_frame_line_pixel_0_0_4 = pixelOut_payload_frame_line_pixel_0_0_4;
  assign videoOut_payload_frame_line_pixel_0_0_5 = pixelOut_payload_frame_line_pixel_0_0_5;
  assign videoOut_payload_frame_line_pixel_0_0_6 = pixelOut_payload_frame_line_pixel_0_0_6;
  assign videoOut_payload_frame_line_pixel_0_0_7 = pixelOut_payload_frame_line_pixel_0_0_7;
  assign videoOut_payload_frame_line_pixel_0_0_8 = pixelOut_payload_frame_line_pixel_0_0_8;
  assign videoOut_payload_frame_line_pixel_0_0_9 = pixelOut_payload_frame_line_pixel_0_0_9;
  assign videoOut_payload_frame_line_pixel_0_0_10 = pixelOut_payload_frame_line_pixel_0_0_10;
  assign videoOut_payload_frame_line_pixel_0_0_11 = pixelOut_payload_frame_line_pixel_0_0_11;
  assign videoOut_payload_frame_line_pixel_0_0_12 = pixelOut_payload_frame_line_pixel_0_0_12;
  assign videoOut_payload_frame_line_pixel_0_0_13 = pixelOut_payload_frame_line_pixel_0_0_13;
  assign videoOut_payload_frame_line_pixel_0_0_14 = pixelOut_payload_frame_line_pixel_0_0_14;
  assign videoOut_payload_frame_line_pixel_0_0_15 = pixelOut_payload_frame_line_pixel_0_0_15;
  assign videoOut_payload_frame_line_pixel_0_1_0 = pixelOut_payload_frame_line_pixel_1_0_0;
  assign videoOut_payload_frame_line_pixel_0_1_1 = pixelOut_payload_frame_line_pixel_1_0_1;
  assign videoOut_payload_frame_line_pixel_0_1_2 = pixelOut_payload_frame_line_pixel_1_0_2;
  assign videoOut_payload_frame_line_pixel_0_1_3 = pixelOut_payload_frame_line_pixel_1_0_3;
  assign videoOut_payload_frame_line_pixel_0_1_4 = pixelOut_payload_frame_line_pixel_1_0_4;
  assign videoOut_payload_frame_line_pixel_0_1_5 = pixelOut_payload_frame_line_pixel_1_0_5;
  assign videoOut_payload_frame_line_pixel_0_1_6 = pixelOut_payload_frame_line_pixel_1_0_6;
  assign videoOut_payload_frame_line_pixel_0_1_7 = pixelOut_payload_frame_line_pixel_1_0_7;
  assign videoOut_payload_frame_line_pixel_0_1_8 = pixelOut_payload_frame_line_pixel_1_0_8;
  assign videoOut_payload_frame_line_pixel_0_1_9 = pixelOut_payload_frame_line_pixel_1_0_9;
  assign videoOut_payload_frame_line_pixel_0_1_10 = pixelOut_payload_frame_line_pixel_1_0_10;
  assign videoOut_payload_frame_line_pixel_0_1_11 = pixelOut_payload_frame_line_pixel_1_0_11;
  assign videoOut_payload_frame_line_pixel_0_1_12 = pixelOut_payload_frame_line_pixel_1_0_12;
  assign videoOut_payload_frame_line_pixel_0_1_13 = pixelOut_payload_frame_line_pixel_1_0_13;
  assign videoOut_payload_frame_line_pixel_0_1_14 = pixelOut_payload_frame_line_pixel_1_0_14;
  assign videoOut_payload_frame_line_pixel_0_1_15 = pixelOut_payload_frame_line_pixel_1_0_15;
  assign videoOut_payload_frame_line_pixel_0_2_0 = pixelOut_payload_frame_line_pixel_2_0_0;
  assign videoOut_payload_frame_line_pixel_0_2_1 = pixelOut_payload_frame_line_pixel_2_0_1;
  assign videoOut_payload_frame_line_pixel_0_2_2 = pixelOut_payload_frame_line_pixel_2_0_2;
  assign videoOut_payload_frame_line_pixel_0_2_3 = pixelOut_payload_frame_line_pixel_2_0_3;
  assign videoOut_payload_frame_line_pixel_0_2_4 = pixelOut_payload_frame_line_pixel_2_0_4;
  assign videoOut_payload_frame_line_pixel_0_2_5 = pixelOut_payload_frame_line_pixel_2_0_5;
  assign videoOut_payload_frame_line_pixel_0_2_6 = pixelOut_payload_frame_line_pixel_2_0_6;
  assign videoOut_payload_frame_line_pixel_0_2_7 = pixelOut_payload_frame_line_pixel_2_0_7;
  assign videoOut_payload_frame_line_pixel_0_2_8 = pixelOut_payload_frame_line_pixel_2_0_8;
  assign videoOut_payload_frame_line_pixel_0_2_9 = pixelOut_payload_frame_line_pixel_2_0_9;
  assign videoOut_payload_frame_line_pixel_0_2_10 = pixelOut_payload_frame_line_pixel_2_0_10;
  assign videoOut_payload_frame_line_pixel_0_2_11 = pixelOut_payload_frame_line_pixel_2_0_11;
  assign videoOut_payload_frame_line_pixel_0_2_12 = pixelOut_payload_frame_line_pixel_2_0_12;
  assign videoOut_payload_frame_line_pixel_0_2_13 = pixelOut_payload_frame_line_pixel_2_0_13;
  assign videoOut_payload_frame_line_pixel_0_2_14 = pixelOut_payload_frame_line_pixel_2_0_14;
  assign videoOut_payload_frame_line_pixel_0_2_15 = pixelOut_payload_frame_line_pixel_2_0_15;
  assign videoOut_payload_frame_line_pixel_1_0_0 = pixelOut_payload_frame_line_pixel_0_1_0;
  assign videoOut_payload_frame_line_pixel_1_0_1 = pixelOut_payload_frame_line_pixel_0_1_1;
  assign videoOut_payload_frame_line_pixel_1_0_2 = pixelOut_payload_frame_line_pixel_0_1_2;
  assign videoOut_payload_frame_line_pixel_1_0_3 = pixelOut_payload_frame_line_pixel_0_1_3;
  assign videoOut_payload_frame_line_pixel_1_0_4 = pixelOut_payload_frame_line_pixel_0_1_4;
  assign videoOut_payload_frame_line_pixel_1_0_5 = pixelOut_payload_frame_line_pixel_0_1_5;
  assign videoOut_payload_frame_line_pixel_1_0_6 = pixelOut_payload_frame_line_pixel_0_1_6;
  assign videoOut_payload_frame_line_pixel_1_0_7 = pixelOut_payload_frame_line_pixel_0_1_7;
  assign videoOut_payload_frame_line_pixel_1_0_8 = pixelOut_payload_frame_line_pixel_0_1_8;
  assign videoOut_payload_frame_line_pixel_1_0_9 = pixelOut_payload_frame_line_pixel_0_1_9;
  assign videoOut_payload_frame_line_pixel_1_0_10 = pixelOut_payload_frame_line_pixel_0_1_10;
  assign videoOut_payload_frame_line_pixel_1_0_11 = pixelOut_payload_frame_line_pixel_0_1_11;
  assign videoOut_payload_frame_line_pixel_1_0_12 = pixelOut_payload_frame_line_pixel_0_1_12;
  assign videoOut_payload_frame_line_pixel_1_0_13 = pixelOut_payload_frame_line_pixel_0_1_13;
  assign videoOut_payload_frame_line_pixel_1_0_14 = pixelOut_payload_frame_line_pixel_0_1_14;
  assign videoOut_payload_frame_line_pixel_1_0_15 = pixelOut_payload_frame_line_pixel_0_1_15;
  assign videoOut_payload_frame_line_pixel_1_1_0 = pixelOut_payload_frame_line_pixel_1_1_0;
  assign videoOut_payload_frame_line_pixel_1_1_1 = pixelOut_payload_frame_line_pixel_1_1_1;
  assign videoOut_payload_frame_line_pixel_1_1_2 = pixelOut_payload_frame_line_pixel_1_1_2;
  assign videoOut_payload_frame_line_pixel_1_1_3 = pixelOut_payload_frame_line_pixel_1_1_3;
  assign videoOut_payload_frame_line_pixel_1_1_4 = pixelOut_payload_frame_line_pixel_1_1_4;
  assign videoOut_payload_frame_line_pixel_1_1_5 = pixelOut_payload_frame_line_pixel_1_1_5;
  assign videoOut_payload_frame_line_pixel_1_1_6 = pixelOut_payload_frame_line_pixel_1_1_6;
  assign videoOut_payload_frame_line_pixel_1_1_7 = pixelOut_payload_frame_line_pixel_1_1_7;
  assign videoOut_payload_frame_line_pixel_1_1_8 = pixelOut_payload_frame_line_pixel_1_1_8;
  assign videoOut_payload_frame_line_pixel_1_1_9 = pixelOut_payload_frame_line_pixel_1_1_9;
  assign videoOut_payload_frame_line_pixel_1_1_10 = pixelOut_payload_frame_line_pixel_1_1_10;
  assign videoOut_payload_frame_line_pixel_1_1_11 = pixelOut_payload_frame_line_pixel_1_1_11;
  assign videoOut_payload_frame_line_pixel_1_1_12 = pixelOut_payload_frame_line_pixel_1_1_12;
  assign videoOut_payload_frame_line_pixel_1_1_13 = pixelOut_payload_frame_line_pixel_1_1_13;
  assign videoOut_payload_frame_line_pixel_1_1_14 = pixelOut_payload_frame_line_pixel_1_1_14;
  assign videoOut_payload_frame_line_pixel_1_1_15 = pixelOut_payload_frame_line_pixel_1_1_15;
  assign videoOut_payload_frame_line_pixel_1_2_0 = pixelOut_payload_frame_line_pixel_2_1_0;
  assign videoOut_payload_frame_line_pixel_1_2_1 = pixelOut_payload_frame_line_pixel_2_1_1;
  assign videoOut_payload_frame_line_pixel_1_2_2 = pixelOut_payload_frame_line_pixel_2_1_2;
  assign videoOut_payload_frame_line_pixel_1_2_3 = pixelOut_payload_frame_line_pixel_2_1_3;
  assign videoOut_payload_frame_line_pixel_1_2_4 = pixelOut_payload_frame_line_pixel_2_1_4;
  assign videoOut_payload_frame_line_pixel_1_2_5 = pixelOut_payload_frame_line_pixel_2_1_5;
  assign videoOut_payload_frame_line_pixel_1_2_6 = pixelOut_payload_frame_line_pixel_2_1_6;
  assign videoOut_payload_frame_line_pixel_1_2_7 = pixelOut_payload_frame_line_pixel_2_1_7;
  assign videoOut_payload_frame_line_pixel_1_2_8 = pixelOut_payload_frame_line_pixel_2_1_8;
  assign videoOut_payload_frame_line_pixel_1_2_9 = pixelOut_payload_frame_line_pixel_2_1_9;
  assign videoOut_payload_frame_line_pixel_1_2_10 = pixelOut_payload_frame_line_pixel_2_1_10;
  assign videoOut_payload_frame_line_pixel_1_2_11 = pixelOut_payload_frame_line_pixel_2_1_11;
  assign videoOut_payload_frame_line_pixel_1_2_12 = pixelOut_payload_frame_line_pixel_2_1_12;
  assign videoOut_payload_frame_line_pixel_1_2_13 = pixelOut_payload_frame_line_pixel_2_1_13;
  assign videoOut_payload_frame_line_pixel_1_2_14 = pixelOut_payload_frame_line_pixel_2_1_14;
  assign videoOut_payload_frame_line_pixel_1_2_15 = pixelOut_payload_frame_line_pixel_2_1_15;
  assign videoOut_payload_frame_line_pixel_2_0_0 = pixelOut_payload_frame_line_pixel_0_2_0;
  assign videoOut_payload_frame_line_pixel_2_0_1 = pixelOut_payload_frame_line_pixel_0_2_1;
  assign videoOut_payload_frame_line_pixel_2_0_2 = pixelOut_payload_frame_line_pixel_0_2_2;
  assign videoOut_payload_frame_line_pixel_2_0_3 = pixelOut_payload_frame_line_pixel_0_2_3;
  assign videoOut_payload_frame_line_pixel_2_0_4 = pixelOut_payload_frame_line_pixel_0_2_4;
  assign videoOut_payload_frame_line_pixel_2_0_5 = pixelOut_payload_frame_line_pixel_0_2_5;
  assign videoOut_payload_frame_line_pixel_2_0_6 = pixelOut_payload_frame_line_pixel_0_2_6;
  assign videoOut_payload_frame_line_pixel_2_0_7 = pixelOut_payload_frame_line_pixel_0_2_7;
  assign videoOut_payload_frame_line_pixel_2_0_8 = pixelOut_payload_frame_line_pixel_0_2_8;
  assign videoOut_payload_frame_line_pixel_2_0_9 = pixelOut_payload_frame_line_pixel_0_2_9;
  assign videoOut_payload_frame_line_pixel_2_0_10 = pixelOut_payload_frame_line_pixel_0_2_10;
  assign videoOut_payload_frame_line_pixel_2_0_11 = pixelOut_payload_frame_line_pixel_0_2_11;
  assign videoOut_payload_frame_line_pixel_2_0_12 = pixelOut_payload_frame_line_pixel_0_2_12;
  assign videoOut_payload_frame_line_pixel_2_0_13 = pixelOut_payload_frame_line_pixel_0_2_13;
  assign videoOut_payload_frame_line_pixel_2_0_14 = pixelOut_payload_frame_line_pixel_0_2_14;
  assign videoOut_payload_frame_line_pixel_2_0_15 = pixelOut_payload_frame_line_pixel_0_2_15;
  assign videoOut_payload_frame_line_pixel_2_1_0 = pixelOut_payload_frame_line_pixel_1_2_0;
  assign videoOut_payload_frame_line_pixel_2_1_1 = pixelOut_payload_frame_line_pixel_1_2_1;
  assign videoOut_payload_frame_line_pixel_2_1_2 = pixelOut_payload_frame_line_pixel_1_2_2;
  assign videoOut_payload_frame_line_pixel_2_1_3 = pixelOut_payload_frame_line_pixel_1_2_3;
  assign videoOut_payload_frame_line_pixel_2_1_4 = pixelOut_payload_frame_line_pixel_1_2_4;
  assign videoOut_payload_frame_line_pixel_2_1_5 = pixelOut_payload_frame_line_pixel_1_2_5;
  assign videoOut_payload_frame_line_pixel_2_1_6 = pixelOut_payload_frame_line_pixel_1_2_6;
  assign videoOut_payload_frame_line_pixel_2_1_7 = pixelOut_payload_frame_line_pixel_1_2_7;
  assign videoOut_payload_frame_line_pixel_2_1_8 = pixelOut_payload_frame_line_pixel_1_2_8;
  assign videoOut_payload_frame_line_pixel_2_1_9 = pixelOut_payload_frame_line_pixel_1_2_9;
  assign videoOut_payload_frame_line_pixel_2_1_10 = pixelOut_payload_frame_line_pixel_1_2_10;
  assign videoOut_payload_frame_line_pixel_2_1_11 = pixelOut_payload_frame_line_pixel_1_2_11;
  assign videoOut_payload_frame_line_pixel_2_1_12 = pixelOut_payload_frame_line_pixel_1_2_12;
  assign videoOut_payload_frame_line_pixel_2_1_13 = pixelOut_payload_frame_line_pixel_1_2_13;
  assign videoOut_payload_frame_line_pixel_2_1_14 = pixelOut_payload_frame_line_pixel_1_2_14;
  assign videoOut_payload_frame_line_pixel_2_1_15 = pixelOut_payload_frame_line_pixel_1_2_15;
  assign videoOut_payload_frame_line_pixel_2_2_0 = pixelOut_payload_frame_line_pixel_2_2_0;
  assign videoOut_payload_frame_line_pixel_2_2_1 = pixelOut_payload_frame_line_pixel_2_2_1;
  assign videoOut_payload_frame_line_pixel_2_2_2 = pixelOut_payload_frame_line_pixel_2_2_2;
  assign videoOut_payload_frame_line_pixel_2_2_3 = pixelOut_payload_frame_line_pixel_2_2_3;
  assign videoOut_payload_frame_line_pixel_2_2_4 = pixelOut_payload_frame_line_pixel_2_2_4;
  assign videoOut_payload_frame_line_pixel_2_2_5 = pixelOut_payload_frame_line_pixel_2_2_5;
  assign videoOut_payload_frame_line_pixel_2_2_6 = pixelOut_payload_frame_line_pixel_2_2_6;
  assign videoOut_payload_frame_line_pixel_2_2_7 = pixelOut_payload_frame_line_pixel_2_2_7;
  assign videoOut_payload_frame_line_pixel_2_2_8 = pixelOut_payload_frame_line_pixel_2_2_8;
  assign videoOut_payload_frame_line_pixel_2_2_9 = pixelOut_payload_frame_line_pixel_2_2_9;
  assign videoOut_payload_frame_line_pixel_2_2_10 = pixelOut_payload_frame_line_pixel_2_2_10;
  assign videoOut_payload_frame_line_pixel_2_2_11 = pixelOut_payload_frame_line_pixel_2_2_11;
  assign videoOut_payload_frame_line_pixel_2_2_12 = pixelOut_payload_frame_line_pixel_2_2_12;
  assign videoOut_payload_frame_line_pixel_2_2_13 = pixelOut_payload_frame_line_pixel_2_2_13;
  assign videoOut_payload_frame_line_pixel_2_2_14 = pixelOut_payload_frame_line_pixel_2_2_14;
  assign videoOut_payload_frame_line_pixel_2_2_15 = pixelOut_payload_frame_line_pixel_2_2_15;
  always @(posedge clk) begin
    if(reset) begin
      pixel_videoOut_rValid <= 1'b0;
      line_videoOut_rValid <= 1'b0;
      line_videoOut_m2sPipe_rValid <= 1'b0;
    end else begin
      if(pixel_videoOut_ready) begin
        pixel_videoOut_rValid <= pixel_videoOut_valid;
      end
      if(line_videoOut_ready) begin
        line_videoOut_rValid <= line_videoOut_valid;
      end
      if(line_videoOut_m2sPipe_valid) begin
        line_videoOut_m2sPipe_rValid <= 1'b1;
      end
      if(line_videoOut_m2sPipe_s2mPipe_ready) begin
        line_videoOut_m2sPipe_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(pixel_videoOut_ready) begin
      pixel_videoOut_rData_frame_line_pixel_0_0_0 <= pixel_videoOut_payload_frame_line_pixel_0_0_0;
      pixel_videoOut_rData_frame_line_pixel_0_0_1 <= pixel_videoOut_payload_frame_line_pixel_0_0_1;
      pixel_videoOut_rData_frame_line_pixel_0_0_2 <= pixel_videoOut_payload_frame_line_pixel_0_0_2;
      pixel_videoOut_rData_frame_line_pixel_0_0_3 <= pixel_videoOut_payload_frame_line_pixel_0_0_3;
      pixel_videoOut_rData_frame_line_pixel_0_0_4 <= pixel_videoOut_payload_frame_line_pixel_0_0_4;
      pixel_videoOut_rData_frame_line_pixel_0_0_5 <= pixel_videoOut_payload_frame_line_pixel_0_0_5;
      pixel_videoOut_rData_frame_line_pixel_0_0_6 <= pixel_videoOut_payload_frame_line_pixel_0_0_6;
      pixel_videoOut_rData_frame_line_pixel_0_0_7 <= pixel_videoOut_payload_frame_line_pixel_0_0_7;
      pixel_videoOut_rData_frame_line_pixel_0_0_8 <= pixel_videoOut_payload_frame_line_pixel_0_0_8;
      pixel_videoOut_rData_frame_line_pixel_0_0_9 <= pixel_videoOut_payload_frame_line_pixel_0_0_9;
      pixel_videoOut_rData_frame_line_pixel_0_0_10 <= pixel_videoOut_payload_frame_line_pixel_0_0_10;
      pixel_videoOut_rData_frame_line_pixel_0_0_11 <= pixel_videoOut_payload_frame_line_pixel_0_0_11;
      pixel_videoOut_rData_frame_line_pixel_0_0_12 <= pixel_videoOut_payload_frame_line_pixel_0_0_12;
      pixel_videoOut_rData_frame_line_pixel_0_0_13 <= pixel_videoOut_payload_frame_line_pixel_0_0_13;
      pixel_videoOut_rData_frame_line_pixel_0_0_14 <= pixel_videoOut_payload_frame_line_pixel_0_0_14;
      pixel_videoOut_rData_frame_line_pixel_0_0_15 <= pixel_videoOut_payload_frame_line_pixel_0_0_15;
      pixel_videoOut_rData_frame_line_pixel_0_1_0 <= pixel_videoOut_payload_frame_line_pixel_0_1_0;
      pixel_videoOut_rData_frame_line_pixel_0_1_1 <= pixel_videoOut_payload_frame_line_pixel_0_1_1;
      pixel_videoOut_rData_frame_line_pixel_0_1_2 <= pixel_videoOut_payload_frame_line_pixel_0_1_2;
      pixel_videoOut_rData_frame_line_pixel_0_1_3 <= pixel_videoOut_payload_frame_line_pixel_0_1_3;
      pixel_videoOut_rData_frame_line_pixel_0_1_4 <= pixel_videoOut_payload_frame_line_pixel_0_1_4;
      pixel_videoOut_rData_frame_line_pixel_0_1_5 <= pixel_videoOut_payload_frame_line_pixel_0_1_5;
      pixel_videoOut_rData_frame_line_pixel_0_1_6 <= pixel_videoOut_payload_frame_line_pixel_0_1_6;
      pixel_videoOut_rData_frame_line_pixel_0_1_7 <= pixel_videoOut_payload_frame_line_pixel_0_1_7;
      pixel_videoOut_rData_frame_line_pixel_0_1_8 <= pixel_videoOut_payload_frame_line_pixel_0_1_8;
      pixel_videoOut_rData_frame_line_pixel_0_1_9 <= pixel_videoOut_payload_frame_line_pixel_0_1_9;
      pixel_videoOut_rData_frame_line_pixel_0_1_10 <= pixel_videoOut_payload_frame_line_pixel_0_1_10;
      pixel_videoOut_rData_frame_line_pixel_0_1_11 <= pixel_videoOut_payload_frame_line_pixel_0_1_11;
      pixel_videoOut_rData_frame_line_pixel_0_1_12 <= pixel_videoOut_payload_frame_line_pixel_0_1_12;
      pixel_videoOut_rData_frame_line_pixel_0_1_13 <= pixel_videoOut_payload_frame_line_pixel_0_1_13;
      pixel_videoOut_rData_frame_line_pixel_0_1_14 <= pixel_videoOut_payload_frame_line_pixel_0_1_14;
      pixel_videoOut_rData_frame_line_pixel_0_1_15 <= pixel_videoOut_payload_frame_line_pixel_0_1_15;
      pixel_videoOut_rData_frame_line_pixel_0_2_0 <= pixel_videoOut_payload_frame_line_pixel_0_2_0;
      pixel_videoOut_rData_frame_line_pixel_0_2_1 <= pixel_videoOut_payload_frame_line_pixel_0_2_1;
      pixel_videoOut_rData_frame_line_pixel_0_2_2 <= pixel_videoOut_payload_frame_line_pixel_0_2_2;
      pixel_videoOut_rData_frame_line_pixel_0_2_3 <= pixel_videoOut_payload_frame_line_pixel_0_2_3;
      pixel_videoOut_rData_frame_line_pixel_0_2_4 <= pixel_videoOut_payload_frame_line_pixel_0_2_4;
      pixel_videoOut_rData_frame_line_pixel_0_2_5 <= pixel_videoOut_payload_frame_line_pixel_0_2_5;
      pixel_videoOut_rData_frame_line_pixel_0_2_6 <= pixel_videoOut_payload_frame_line_pixel_0_2_6;
      pixel_videoOut_rData_frame_line_pixel_0_2_7 <= pixel_videoOut_payload_frame_line_pixel_0_2_7;
      pixel_videoOut_rData_frame_line_pixel_0_2_8 <= pixel_videoOut_payload_frame_line_pixel_0_2_8;
      pixel_videoOut_rData_frame_line_pixel_0_2_9 <= pixel_videoOut_payload_frame_line_pixel_0_2_9;
      pixel_videoOut_rData_frame_line_pixel_0_2_10 <= pixel_videoOut_payload_frame_line_pixel_0_2_10;
      pixel_videoOut_rData_frame_line_pixel_0_2_11 <= pixel_videoOut_payload_frame_line_pixel_0_2_11;
      pixel_videoOut_rData_frame_line_pixel_0_2_12 <= pixel_videoOut_payload_frame_line_pixel_0_2_12;
      pixel_videoOut_rData_frame_line_pixel_0_2_13 <= pixel_videoOut_payload_frame_line_pixel_0_2_13;
      pixel_videoOut_rData_frame_line_pixel_0_2_14 <= pixel_videoOut_payload_frame_line_pixel_0_2_14;
      pixel_videoOut_rData_frame_line_pixel_0_2_15 <= pixel_videoOut_payload_frame_line_pixel_0_2_15;
      pixel_videoOut_rData_frame_line_pixel_1_0_0 <= pixel_videoOut_payload_frame_line_pixel_1_0_0;
      pixel_videoOut_rData_frame_line_pixel_1_0_1 <= pixel_videoOut_payload_frame_line_pixel_1_0_1;
      pixel_videoOut_rData_frame_line_pixel_1_0_2 <= pixel_videoOut_payload_frame_line_pixel_1_0_2;
      pixel_videoOut_rData_frame_line_pixel_1_0_3 <= pixel_videoOut_payload_frame_line_pixel_1_0_3;
      pixel_videoOut_rData_frame_line_pixel_1_0_4 <= pixel_videoOut_payload_frame_line_pixel_1_0_4;
      pixel_videoOut_rData_frame_line_pixel_1_0_5 <= pixel_videoOut_payload_frame_line_pixel_1_0_5;
      pixel_videoOut_rData_frame_line_pixel_1_0_6 <= pixel_videoOut_payload_frame_line_pixel_1_0_6;
      pixel_videoOut_rData_frame_line_pixel_1_0_7 <= pixel_videoOut_payload_frame_line_pixel_1_0_7;
      pixel_videoOut_rData_frame_line_pixel_1_0_8 <= pixel_videoOut_payload_frame_line_pixel_1_0_8;
      pixel_videoOut_rData_frame_line_pixel_1_0_9 <= pixel_videoOut_payload_frame_line_pixel_1_0_9;
      pixel_videoOut_rData_frame_line_pixel_1_0_10 <= pixel_videoOut_payload_frame_line_pixel_1_0_10;
      pixel_videoOut_rData_frame_line_pixel_1_0_11 <= pixel_videoOut_payload_frame_line_pixel_1_0_11;
      pixel_videoOut_rData_frame_line_pixel_1_0_12 <= pixel_videoOut_payload_frame_line_pixel_1_0_12;
      pixel_videoOut_rData_frame_line_pixel_1_0_13 <= pixel_videoOut_payload_frame_line_pixel_1_0_13;
      pixel_videoOut_rData_frame_line_pixel_1_0_14 <= pixel_videoOut_payload_frame_line_pixel_1_0_14;
      pixel_videoOut_rData_frame_line_pixel_1_0_15 <= pixel_videoOut_payload_frame_line_pixel_1_0_15;
      pixel_videoOut_rData_frame_line_pixel_1_1_0 <= pixel_videoOut_payload_frame_line_pixel_1_1_0;
      pixel_videoOut_rData_frame_line_pixel_1_1_1 <= pixel_videoOut_payload_frame_line_pixel_1_1_1;
      pixel_videoOut_rData_frame_line_pixel_1_1_2 <= pixel_videoOut_payload_frame_line_pixel_1_1_2;
      pixel_videoOut_rData_frame_line_pixel_1_1_3 <= pixel_videoOut_payload_frame_line_pixel_1_1_3;
      pixel_videoOut_rData_frame_line_pixel_1_1_4 <= pixel_videoOut_payload_frame_line_pixel_1_1_4;
      pixel_videoOut_rData_frame_line_pixel_1_1_5 <= pixel_videoOut_payload_frame_line_pixel_1_1_5;
      pixel_videoOut_rData_frame_line_pixel_1_1_6 <= pixel_videoOut_payload_frame_line_pixel_1_1_6;
      pixel_videoOut_rData_frame_line_pixel_1_1_7 <= pixel_videoOut_payload_frame_line_pixel_1_1_7;
      pixel_videoOut_rData_frame_line_pixel_1_1_8 <= pixel_videoOut_payload_frame_line_pixel_1_1_8;
      pixel_videoOut_rData_frame_line_pixel_1_1_9 <= pixel_videoOut_payload_frame_line_pixel_1_1_9;
      pixel_videoOut_rData_frame_line_pixel_1_1_10 <= pixel_videoOut_payload_frame_line_pixel_1_1_10;
      pixel_videoOut_rData_frame_line_pixel_1_1_11 <= pixel_videoOut_payload_frame_line_pixel_1_1_11;
      pixel_videoOut_rData_frame_line_pixel_1_1_12 <= pixel_videoOut_payload_frame_line_pixel_1_1_12;
      pixel_videoOut_rData_frame_line_pixel_1_1_13 <= pixel_videoOut_payload_frame_line_pixel_1_1_13;
      pixel_videoOut_rData_frame_line_pixel_1_1_14 <= pixel_videoOut_payload_frame_line_pixel_1_1_14;
      pixel_videoOut_rData_frame_line_pixel_1_1_15 <= pixel_videoOut_payload_frame_line_pixel_1_1_15;
      pixel_videoOut_rData_frame_line_pixel_1_2_0 <= pixel_videoOut_payload_frame_line_pixel_1_2_0;
      pixel_videoOut_rData_frame_line_pixel_1_2_1 <= pixel_videoOut_payload_frame_line_pixel_1_2_1;
      pixel_videoOut_rData_frame_line_pixel_1_2_2 <= pixel_videoOut_payload_frame_line_pixel_1_2_2;
      pixel_videoOut_rData_frame_line_pixel_1_2_3 <= pixel_videoOut_payload_frame_line_pixel_1_2_3;
      pixel_videoOut_rData_frame_line_pixel_1_2_4 <= pixel_videoOut_payload_frame_line_pixel_1_2_4;
      pixel_videoOut_rData_frame_line_pixel_1_2_5 <= pixel_videoOut_payload_frame_line_pixel_1_2_5;
      pixel_videoOut_rData_frame_line_pixel_1_2_6 <= pixel_videoOut_payload_frame_line_pixel_1_2_6;
      pixel_videoOut_rData_frame_line_pixel_1_2_7 <= pixel_videoOut_payload_frame_line_pixel_1_2_7;
      pixel_videoOut_rData_frame_line_pixel_1_2_8 <= pixel_videoOut_payload_frame_line_pixel_1_2_8;
      pixel_videoOut_rData_frame_line_pixel_1_2_9 <= pixel_videoOut_payload_frame_line_pixel_1_2_9;
      pixel_videoOut_rData_frame_line_pixel_1_2_10 <= pixel_videoOut_payload_frame_line_pixel_1_2_10;
      pixel_videoOut_rData_frame_line_pixel_1_2_11 <= pixel_videoOut_payload_frame_line_pixel_1_2_11;
      pixel_videoOut_rData_frame_line_pixel_1_2_12 <= pixel_videoOut_payload_frame_line_pixel_1_2_12;
      pixel_videoOut_rData_frame_line_pixel_1_2_13 <= pixel_videoOut_payload_frame_line_pixel_1_2_13;
      pixel_videoOut_rData_frame_line_pixel_1_2_14 <= pixel_videoOut_payload_frame_line_pixel_1_2_14;
      pixel_videoOut_rData_frame_line_pixel_1_2_15 <= pixel_videoOut_payload_frame_line_pixel_1_2_15;
      pixel_videoOut_rData_frame_line_pixel_2_0_0 <= pixel_videoOut_payload_frame_line_pixel_2_0_0;
      pixel_videoOut_rData_frame_line_pixel_2_0_1 <= pixel_videoOut_payload_frame_line_pixel_2_0_1;
      pixel_videoOut_rData_frame_line_pixel_2_0_2 <= pixel_videoOut_payload_frame_line_pixel_2_0_2;
      pixel_videoOut_rData_frame_line_pixel_2_0_3 <= pixel_videoOut_payload_frame_line_pixel_2_0_3;
      pixel_videoOut_rData_frame_line_pixel_2_0_4 <= pixel_videoOut_payload_frame_line_pixel_2_0_4;
      pixel_videoOut_rData_frame_line_pixel_2_0_5 <= pixel_videoOut_payload_frame_line_pixel_2_0_5;
      pixel_videoOut_rData_frame_line_pixel_2_0_6 <= pixel_videoOut_payload_frame_line_pixel_2_0_6;
      pixel_videoOut_rData_frame_line_pixel_2_0_7 <= pixel_videoOut_payload_frame_line_pixel_2_0_7;
      pixel_videoOut_rData_frame_line_pixel_2_0_8 <= pixel_videoOut_payload_frame_line_pixel_2_0_8;
      pixel_videoOut_rData_frame_line_pixel_2_0_9 <= pixel_videoOut_payload_frame_line_pixel_2_0_9;
      pixel_videoOut_rData_frame_line_pixel_2_0_10 <= pixel_videoOut_payload_frame_line_pixel_2_0_10;
      pixel_videoOut_rData_frame_line_pixel_2_0_11 <= pixel_videoOut_payload_frame_line_pixel_2_0_11;
      pixel_videoOut_rData_frame_line_pixel_2_0_12 <= pixel_videoOut_payload_frame_line_pixel_2_0_12;
      pixel_videoOut_rData_frame_line_pixel_2_0_13 <= pixel_videoOut_payload_frame_line_pixel_2_0_13;
      pixel_videoOut_rData_frame_line_pixel_2_0_14 <= pixel_videoOut_payload_frame_line_pixel_2_0_14;
      pixel_videoOut_rData_frame_line_pixel_2_0_15 <= pixel_videoOut_payload_frame_line_pixel_2_0_15;
      pixel_videoOut_rData_frame_line_pixel_2_1_0 <= pixel_videoOut_payload_frame_line_pixel_2_1_0;
      pixel_videoOut_rData_frame_line_pixel_2_1_1 <= pixel_videoOut_payload_frame_line_pixel_2_1_1;
      pixel_videoOut_rData_frame_line_pixel_2_1_2 <= pixel_videoOut_payload_frame_line_pixel_2_1_2;
      pixel_videoOut_rData_frame_line_pixel_2_1_3 <= pixel_videoOut_payload_frame_line_pixel_2_1_3;
      pixel_videoOut_rData_frame_line_pixel_2_1_4 <= pixel_videoOut_payload_frame_line_pixel_2_1_4;
      pixel_videoOut_rData_frame_line_pixel_2_1_5 <= pixel_videoOut_payload_frame_line_pixel_2_1_5;
      pixel_videoOut_rData_frame_line_pixel_2_1_6 <= pixel_videoOut_payload_frame_line_pixel_2_1_6;
      pixel_videoOut_rData_frame_line_pixel_2_1_7 <= pixel_videoOut_payload_frame_line_pixel_2_1_7;
      pixel_videoOut_rData_frame_line_pixel_2_1_8 <= pixel_videoOut_payload_frame_line_pixel_2_1_8;
      pixel_videoOut_rData_frame_line_pixel_2_1_9 <= pixel_videoOut_payload_frame_line_pixel_2_1_9;
      pixel_videoOut_rData_frame_line_pixel_2_1_10 <= pixel_videoOut_payload_frame_line_pixel_2_1_10;
      pixel_videoOut_rData_frame_line_pixel_2_1_11 <= pixel_videoOut_payload_frame_line_pixel_2_1_11;
      pixel_videoOut_rData_frame_line_pixel_2_1_12 <= pixel_videoOut_payload_frame_line_pixel_2_1_12;
      pixel_videoOut_rData_frame_line_pixel_2_1_13 <= pixel_videoOut_payload_frame_line_pixel_2_1_13;
      pixel_videoOut_rData_frame_line_pixel_2_1_14 <= pixel_videoOut_payload_frame_line_pixel_2_1_14;
      pixel_videoOut_rData_frame_line_pixel_2_1_15 <= pixel_videoOut_payload_frame_line_pixel_2_1_15;
      pixel_videoOut_rData_frame_line_pixel_2_2_0 <= pixel_videoOut_payload_frame_line_pixel_2_2_0;
      pixel_videoOut_rData_frame_line_pixel_2_2_1 <= pixel_videoOut_payload_frame_line_pixel_2_2_1;
      pixel_videoOut_rData_frame_line_pixel_2_2_2 <= pixel_videoOut_payload_frame_line_pixel_2_2_2;
      pixel_videoOut_rData_frame_line_pixel_2_2_3 <= pixel_videoOut_payload_frame_line_pixel_2_2_3;
      pixel_videoOut_rData_frame_line_pixel_2_2_4 <= pixel_videoOut_payload_frame_line_pixel_2_2_4;
      pixel_videoOut_rData_frame_line_pixel_2_2_5 <= pixel_videoOut_payload_frame_line_pixel_2_2_5;
      pixel_videoOut_rData_frame_line_pixel_2_2_6 <= pixel_videoOut_payload_frame_line_pixel_2_2_6;
      pixel_videoOut_rData_frame_line_pixel_2_2_7 <= pixel_videoOut_payload_frame_line_pixel_2_2_7;
      pixel_videoOut_rData_frame_line_pixel_2_2_8 <= pixel_videoOut_payload_frame_line_pixel_2_2_8;
      pixel_videoOut_rData_frame_line_pixel_2_2_9 <= pixel_videoOut_payload_frame_line_pixel_2_2_9;
      pixel_videoOut_rData_frame_line_pixel_2_2_10 <= pixel_videoOut_payload_frame_line_pixel_2_2_10;
      pixel_videoOut_rData_frame_line_pixel_2_2_11 <= pixel_videoOut_payload_frame_line_pixel_2_2_11;
      pixel_videoOut_rData_frame_line_pixel_2_2_12 <= pixel_videoOut_payload_frame_line_pixel_2_2_12;
      pixel_videoOut_rData_frame_line_pixel_2_2_13 <= pixel_videoOut_payload_frame_line_pixel_2_2_13;
      pixel_videoOut_rData_frame_line_pixel_2_2_14 <= pixel_videoOut_payload_frame_line_pixel_2_2_14;
      pixel_videoOut_rData_frame_line_pixel_2_2_15 <= pixel_videoOut_payload_frame_line_pixel_2_2_15;
      pixel_videoOut_rData_frame_line_endOfLine <= pixel_videoOut_payload_frame_line_endOfLine;
      pixel_videoOut_rData_frame_endOfFrame <= pixel_videoOut_payload_frame_endOfFrame;
      pixel_videoOut_rData_endOfPack <= pixel_videoOut_payload_endOfPack;
    end
    if(line_videoOut_ready) begin
      line_videoOut_rData_frame_line_pixel_0_0 <= line_videoOut_payload_frame_line_pixel_0_0;
      line_videoOut_rData_frame_line_pixel_0_1 <= line_videoOut_payload_frame_line_pixel_0_1;
      line_videoOut_rData_frame_line_pixel_0_2 <= line_videoOut_payload_frame_line_pixel_0_2;
      line_videoOut_rData_frame_line_pixel_0_3 <= line_videoOut_payload_frame_line_pixel_0_3;
      line_videoOut_rData_frame_line_pixel_0_4 <= line_videoOut_payload_frame_line_pixel_0_4;
      line_videoOut_rData_frame_line_pixel_0_5 <= line_videoOut_payload_frame_line_pixel_0_5;
      line_videoOut_rData_frame_line_pixel_0_6 <= line_videoOut_payload_frame_line_pixel_0_6;
      line_videoOut_rData_frame_line_pixel_0_7 <= line_videoOut_payload_frame_line_pixel_0_7;
      line_videoOut_rData_frame_line_pixel_0_8 <= line_videoOut_payload_frame_line_pixel_0_8;
      line_videoOut_rData_frame_line_pixel_0_9 <= line_videoOut_payload_frame_line_pixel_0_9;
      line_videoOut_rData_frame_line_pixel_0_10 <= line_videoOut_payload_frame_line_pixel_0_10;
      line_videoOut_rData_frame_line_pixel_0_11 <= line_videoOut_payload_frame_line_pixel_0_11;
      line_videoOut_rData_frame_line_pixel_0_12 <= line_videoOut_payload_frame_line_pixel_0_12;
      line_videoOut_rData_frame_line_pixel_0_13 <= line_videoOut_payload_frame_line_pixel_0_13;
      line_videoOut_rData_frame_line_pixel_0_14 <= line_videoOut_payload_frame_line_pixel_0_14;
      line_videoOut_rData_frame_line_pixel_0_15 <= line_videoOut_payload_frame_line_pixel_0_15;
      line_videoOut_rData_frame_line_pixel_1_0 <= line_videoOut_payload_frame_line_pixel_1_0;
      line_videoOut_rData_frame_line_pixel_1_1 <= line_videoOut_payload_frame_line_pixel_1_1;
      line_videoOut_rData_frame_line_pixel_1_2 <= line_videoOut_payload_frame_line_pixel_1_2;
      line_videoOut_rData_frame_line_pixel_1_3 <= line_videoOut_payload_frame_line_pixel_1_3;
      line_videoOut_rData_frame_line_pixel_1_4 <= line_videoOut_payload_frame_line_pixel_1_4;
      line_videoOut_rData_frame_line_pixel_1_5 <= line_videoOut_payload_frame_line_pixel_1_5;
      line_videoOut_rData_frame_line_pixel_1_6 <= line_videoOut_payload_frame_line_pixel_1_6;
      line_videoOut_rData_frame_line_pixel_1_7 <= line_videoOut_payload_frame_line_pixel_1_7;
      line_videoOut_rData_frame_line_pixel_1_8 <= line_videoOut_payload_frame_line_pixel_1_8;
      line_videoOut_rData_frame_line_pixel_1_9 <= line_videoOut_payload_frame_line_pixel_1_9;
      line_videoOut_rData_frame_line_pixel_1_10 <= line_videoOut_payload_frame_line_pixel_1_10;
      line_videoOut_rData_frame_line_pixel_1_11 <= line_videoOut_payload_frame_line_pixel_1_11;
      line_videoOut_rData_frame_line_pixel_1_12 <= line_videoOut_payload_frame_line_pixel_1_12;
      line_videoOut_rData_frame_line_pixel_1_13 <= line_videoOut_payload_frame_line_pixel_1_13;
      line_videoOut_rData_frame_line_pixel_1_14 <= line_videoOut_payload_frame_line_pixel_1_14;
      line_videoOut_rData_frame_line_pixel_1_15 <= line_videoOut_payload_frame_line_pixel_1_15;
      line_videoOut_rData_frame_line_pixel_2_0 <= line_videoOut_payload_frame_line_pixel_2_0;
      line_videoOut_rData_frame_line_pixel_2_1 <= line_videoOut_payload_frame_line_pixel_2_1;
      line_videoOut_rData_frame_line_pixel_2_2 <= line_videoOut_payload_frame_line_pixel_2_2;
      line_videoOut_rData_frame_line_pixel_2_3 <= line_videoOut_payload_frame_line_pixel_2_3;
      line_videoOut_rData_frame_line_pixel_2_4 <= line_videoOut_payload_frame_line_pixel_2_4;
      line_videoOut_rData_frame_line_pixel_2_5 <= line_videoOut_payload_frame_line_pixel_2_5;
      line_videoOut_rData_frame_line_pixel_2_6 <= line_videoOut_payload_frame_line_pixel_2_6;
      line_videoOut_rData_frame_line_pixel_2_7 <= line_videoOut_payload_frame_line_pixel_2_7;
      line_videoOut_rData_frame_line_pixel_2_8 <= line_videoOut_payload_frame_line_pixel_2_8;
      line_videoOut_rData_frame_line_pixel_2_9 <= line_videoOut_payload_frame_line_pixel_2_9;
      line_videoOut_rData_frame_line_pixel_2_10 <= line_videoOut_payload_frame_line_pixel_2_10;
      line_videoOut_rData_frame_line_pixel_2_11 <= line_videoOut_payload_frame_line_pixel_2_11;
      line_videoOut_rData_frame_line_pixel_2_12 <= line_videoOut_payload_frame_line_pixel_2_12;
      line_videoOut_rData_frame_line_pixel_2_13 <= line_videoOut_payload_frame_line_pixel_2_13;
      line_videoOut_rData_frame_line_pixel_2_14 <= line_videoOut_payload_frame_line_pixel_2_14;
      line_videoOut_rData_frame_line_pixel_2_15 <= line_videoOut_payload_frame_line_pixel_2_15;
      line_videoOut_rData_frame_line_endOfLine <= line_videoOut_payload_frame_line_endOfLine;
      line_videoOut_rData_frame_endOfFrame <= line_videoOut_payload_frame_endOfFrame;
      line_videoOut_rData_endOfPack <= line_videoOut_payload_endOfPack;
    end
    if(line_videoOut_m2sPipe_ready) begin
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_0 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_0;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_1 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_1;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_2 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_2;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_3 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_3;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_4 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_4;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_5 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_5;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_6 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_6;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_7 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_7;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_8 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_8;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_9 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_9;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_10 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_10;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_11 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_11;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_12 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_12;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_13 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_13;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_14 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_14;
      line_videoOut_m2sPipe_rData_frame_line_pixel_0_15 <= line_videoOut_m2sPipe_payload_frame_line_pixel_0_15;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_0 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_0;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_1 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_1;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_2 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_2;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_3 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_3;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_4 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_4;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_5 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_5;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_6 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_6;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_7 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_7;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_8 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_8;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_9 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_9;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_10 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_10;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_11 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_11;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_12 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_12;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_13 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_13;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_14 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_14;
      line_videoOut_m2sPipe_rData_frame_line_pixel_1_15 <= line_videoOut_m2sPipe_payload_frame_line_pixel_1_15;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_0 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_0;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_1 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_1;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_2 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_2;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_3 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_3;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_4 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_4;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_5 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_5;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_6 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_6;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_7 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_7;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_8 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_8;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_9 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_9;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_10 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_10;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_11 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_11;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_12 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_12;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_13 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_13;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_14 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_14;
      line_videoOut_m2sPipe_rData_frame_line_pixel_2_15 <= line_videoOut_m2sPipe_payload_frame_line_pixel_2_15;
      line_videoOut_m2sPipe_rData_frame_line_endOfLine <= line_videoOut_m2sPipe_payload_frame_line_endOfLine;
      line_videoOut_m2sPipe_rData_frame_endOfFrame <= line_videoOut_m2sPipe_payload_frame_endOfFrame;
      line_videoOut_m2sPipe_rData_endOfPack <= line_videoOut_m2sPipe_payload_endOfPack;
    end
  end


endmodule

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

//StreamFifoHighPerf_2 replaced by StreamFifoHighPerf_2

module StreamFifoHighPerf_2 (
  input               push_valid,
  output              push_ready,
  input      [7:0]    push_payload_0_0_0_0,
  input      [7:0]    push_payload_0_0_0_1,
  input      [7:0]    push_payload_0_0_0_2,
  input      [7:0]    push_payload_0_0_0_3,
  input      [7:0]    push_payload_0_0_0_4,
  input      [7:0]    push_payload_0_0_0_5,
  input      [7:0]    push_payload_0_0_0_6,
  input      [7:0]    push_payload_0_0_0_7,
  input      [7:0]    push_payload_0_0_0_8,
  input      [7:0]    push_payload_0_0_0_9,
  input      [7:0]    push_payload_0_0_0_10,
  input      [7:0]    push_payload_0_0_0_11,
  input      [7:0]    push_payload_0_0_0_12,
  input      [7:0]    push_payload_0_0_0_13,
  input      [7:0]    push_payload_0_0_0_14,
  input      [7:0]    push_payload_0_0_0_15,
  input      [7:0]    push_payload_0_0_1_0,
  input      [7:0]    push_payload_0_0_1_1,
  input      [7:0]    push_payload_0_0_1_2,
  input      [7:0]    push_payload_0_0_1_3,
  input      [7:0]    push_payload_0_0_1_4,
  input      [7:0]    push_payload_0_0_1_5,
  input      [7:0]    push_payload_0_0_1_6,
  input      [7:0]    push_payload_0_0_1_7,
  input      [7:0]    push_payload_0_0_1_8,
  input      [7:0]    push_payload_0_0_1_9,
  input      [7:0]    push_payload_0_0_1_10,
  input      [7:0]    push_payload_0_0_1_11,
  input      [7:0]    push_payload_0_0_1_12,
  input      [7:0]    push_payload_0_0_1_13,
  input      [7:0]    push_payload_0_0_1_14,
  input      [7:0]    push_payload_0_0_1_15,
  input      [7:0]    push_payload_0_0_2_0,
  input      [7:0]    push_payload_0_0_2_1,
  input      [7:0]    push_payload_0_0_2_2,
  input      [7:0]    push_payload_0_0_2_3,
  input      [7:0]    push_payload_0_0_2_4,
  input      [7:0]    push_payload_0_0_2_5,
  input      [7:0]    push_payload_0_0_2_6,
  input      [7:0]    push_payload_0_0_2_7,
  input      [7:0]    push_payload_0_0_2_8,
  input      [7:0]    push_payload_0_0_2_9,
  input      [7:0]    push_payload_0_0_2_10,
  input      [7:0]    push_payload_0_0_2_11,
  input      [7:0]    push_payload_0_0_2_12,
  input      [7:0]    push_payload_0_0_2_13,
  input      [7:0]    push_payload_0_0_2_14,
  input      [7:0]    push_payload_0_0_2_15,
  input      [7:0]    push_payload_0_1_0_0,
  input      [7:0]    push_payload_0_1_0_1,
  input      [7:0]    push_payload_0_1_0_2,
  input      [7:0]    push_payload_0_1_0_3,
  input      [7:0]    push_payload_0_1_0_4,
  input      [7:0]    push_payload_0_1_0_5,
  input      [7:0]    push_payload_0_1_0_6,
  input      [7:0]    push_payload_0_1_0_7,
  input      [7:0]    push_payload_0_1_0_8,
  input      [7:0]    push_payload_0_1_0_9,
  input      [7:0]    push_payload_0_1_0_10,
  input      [7:0]    push_payload_0_1_0_11,
  input      [7:0]    push_payload_0_1_0_12,
  input      [7:0]    push_payload_0_1_0_13,
  input      [7:0]    push_payload_0_1_0_14,
  input      [7:0]    push_payload_0_1_0_15,
  input      [7:0]    push_payload_0_1_1_0,
  input      [7:0]    push_payload_0_1_1_1,
  input      [7:0]    push_payload_0_1_1_2,
  input      [7:0]    push_payload_0_1_1_3,
  input      [7:0]    push_payload_0_1_1_4,
  input      [7:0]    push_payload_0_1_1_5,
  input      [7:0]    push_payload_0_1_1_6,
  input      [7:0]    push_payload_0_1_1_7,
  input      [7:0]    push_payload_0_1_1_8,
  input      [7:0]    push_payload_0_1_1_9,
  input      [7:0]    push_payload_0_1_1_10,
  input      [7:0]    push_payload_0_1_1_11,
  input      [7:0]    push_payload_0_1_1_12,
  input      [7:0]    push_payload_0_1_1_13,
  input      [7:0]    push_payload_0_1_1_14,
  input      [7:0]    push_payload_0_1_1_15,
  input      [7:0]    push_payload_0_1_2_0,
  input      [7:0]    push_payload_0_1_2_1,
  input      [7:0]    push_payload_0_1_2_2,
  input      [7:0]    push_payload_0_1_2_3,
  input      [7:0]    push_payload_0_1_2_4,
  input      [7:0]    push_payload_0_1_2_5,
  input      [7:0]    push_payload_0_1_2_6,
  input      [7:0]    push_payload_0_1_2_7,
  input      [7:0]    push_payload_0_1_2_8,
  input      [7:0]    push_payload_0_1_2_9,
  input      [7:0]    push_payload_0_1_2_10,
  input      [7:0]    push_payload_0_1_2_11,
  input      [7:0]    push_payload_0_1_2_12,
  input      [7:0]    push_payload_0_1_2_13,
  input      [7:0]    push_payload_0_1_2_14,
  input      [7:0]    push_payload_0_1_2_15,
  input      [7:0]    push_payload_0_2_0_0,
  input      [7:0]    push_payload_0_2_0_1,
  input      [7:0]    push_payload_0_2_0_2,
  input      [7:0]    push_payload_0_2_0_3,
  input      [7:0]    push_payload_0_2_0_4,
  input      [7:0]    push_payload_0_2_0_5,
  input      [7:0]    push_payload_0_2_0_6,
  input      [7:0]    push_payload_0_2_0_7,
  input      [7:0]    push_payload_0_2_0_8,
  input      [7:0]    push_payload_0_2_0_9,
  input      [7:0]    push_payload_0_2_0_10,
  input      [7:0]    push_payload_0_2_0_11,
  input      [7:0]    push_payload_0_2_0_12,
  input      [7:0]    push_payload_0_2_0_13,
  input      [7:0]    push_payload_0_2_0_14,
  input      [7:0]    push_payload_0_2_0_15,
  input      [7:0]    push_payload_0_2_1_0,
  input      [7:0]    push_payload_0_2_1_1,
  input      [7:0]    push_payload_0_2_1_2,
  input      [7:0]    push_payload_0_2_1_3,
  input      [7:0]    push_payload_0_2_1_4,
  input      [7:0]    push_payload_0_2_1_5,
  input      [7:0]    push_payload_0_2_1_6,
  input      [7:0]    push_payload_0_2_1_7,
  input      [7:0]    push_payload_0_2_1_8,
  input      [7:0]    push_payload_0_2_1_9,
  input      [7:0]    push_payload_0_2_1_10,
  input      [7:0]    push_payload_0_2_1_11,
  input      [7:0]    push_payload_0_2_1_12,
  input      [7:0]    push_payload_0_2_1_13,
  input      [7:0]    push_payload_0_2_1_14,
  input      [7:0]    push_payload_0_2_1_15,
  input      [7:0]    push_payload_0_2_2_0,
  input      [7:0]    push_payload_0_2_2_1,
  input      [7:0]    push_payload_0_2_2_2,
  input      [7:0]    push_payload_0_2_2_3,
  input      [7:0]    push_payload_0_2_2_4,
  input      [7:0]    push_payload_0_2_2_5,
  input      [7:0]    push_payload_0_2_2_6,
  input      [7:0]    push_payload_0_2_2_7,
  input      [7:0]    push_payload_0_2_2_8,
  input      [7:0]    push_payload_0_2_2_9,
  input      [7:0]    push_payload_0_2_2_10,
  input      [7:0]    push_payload_0_2_2_11,
  input      [7:0]    push_payload_0_2_2_12,
  input      [7:0]    push_payload_0_2_2_13,
  input      [7:0]    push_payload_0_2_2_14,
  input      [7:0]    push_payload_0_2_2_15,
  input      [7:0]    push_payload_1_0_0_0,
  input      [7:0]    push_payload_1_0_0_1,
  input      [7:0]    push_payload_1_0_0_2,
  input      [7:0]    push_payload_1_0_0_3,
  input      [7:0]    push_payload_1_0_0_4,
  input      [7:0]    push_payload_1_0_0_5,
  input      [7:0]    push_payload_1_0_0_6,
  input      [7:0]    push_payload_1_0_0_7,
  input      [7:0]    push_payload_1_0_0_8,
  input      [7:0]    push_payload_1_0_0_9,
  input      [7:0]    push_payload_1_0_0_10,
  input      [7:0]    push_payload_1_0_0_11,
  input      [7:0]    push_payload_1_0_0_12,
  input      [7:0]    push_payload_1_0_0_13,
  input      [7:0]    push_payload_1_0_0_14,
  input      [7:0]    push_payload_1_0_0_15,
  input      [7:0]    push_payload_1_0_1_0,
  input      [7:0]    push_payload_1_0_1_1,
  input      [7:0]    push_payload_1_0_1_2,
  input      [7:0]    push_payload_1_0_1_3,
  input      [7:0]    push_payload_1_0_1_4,
  input      [7:0]    push_payload_1_0_1_5,
  input      [7:0]    push_payload_1_0_1_6,
  input      [7:0]    push_payload_1_0_1_7,
  input      [7:0]    push_payload_1_0_1_8,
  input      [7:0]    push_payload_1_0_1_9,
  input      [7:0]    push_payload_1_0_1_10,
  input      [7:0]    push_payload_1_0_1_11,
  input      [7:0]    push_payload_1_0_1_12,
  input      [7:0]    push_payload_1_0_1_13,
  input      [7:0]    push_payload_1_0_1_14,
  input      [7:0]    push_payload_1_0_1_15,
  input      [7:0]    push_payload_1_0_2_0,
  input      [7:0]    push_payload_1_0_2_1,
  input      [7:0]    push_payload_1_0_2_2,
  input      [7:0]    push_payload_1_0_2_3,
  input      [7:0]    push_payload_1_0_2_4,
  input      [7:0]    push_payload_1_0_2_5,
  input      [7:0]    push_payload_1_0_2_6,
  input      [7:0]    push_payload_1_0_2_7,
  input      [7:0]    push_payload_1_0_2_8,
  input      [7:0]    push_payload_1_0_2_9,
  input      [7:0]    push_payload_1_0_2_10,
  input      [7:0]    push_payload_1_0_2_11,
  input      [7:0]    push_payload_1_0_2_12,
  input      [7:0]    push_payload_1_0_2_13,
  input      [7:0]    push_payload_1_0_2_14,
  input      [7:0]    push_payload_1_0_2_15,
  input      [7:0]    push_payload_1_1_0_0,
  input      [7:0]    push_payload_1_1_0_1,
  input      [7:0]    push_payload_1_1_0_2,
  input      [7:0]    push_payload_1_1_0_3,
  input      [7:0]    push_payload_1_1_0_4,
  input      [7:0]    push_payload_1_1_0_5,
  input      [7:0]    push_payload_1_1_0_6,
  input      [7:0]    push_payload_1_1_0_7,
  input      [7:0]    push_payload_1_1_0_8,
  input      [7:0]    push_payload_1_1_0_9,
  input      [7:0]    push_payload_1_1_0_10,
  input      [7:0]    push_payload_1_1_0_11,
  input      [7:0]    push_payload_1_1_0_12,
  input      [7:0]    push_payload_1_1_0_13,
  input      [7:0]    push_payload_1_1_0_14,
  input      [7:0]    push_payload_1_1_0_15,
  input      [7:0]    push_payload_1_1_1_0,
  input      [7:0]    push_payload_1_1_1_1,
  input      [7:0]    push_payload_1_1_1_2,
  input      [7:0]    push_payload_1_1_1_3,
  input      [7:0]    push_payload_1_1_1_4,
  input      [7:0]    push_payload_1_1_1_5,
  input      [7:0]    push_payload_1_1_1_6,
  input      [7:0]    push_payload_1_1_1_7,
  input      [7:0]    push_payload_1_1_1_8,
  input      [7:0]    push_payload_1_1_1_9,
  input      [7:0]    push_payload_1_1_1_10,
  input      [7:0]    push_payload_1_1_1_11,
  input      [7:0]    push_payload_1_1_1_12,
  input      [7:0]    push_payload_1_1_1_13,
  input      [7:0]    push_payload_1_1_1_14,
  input      [7:0]    push_payload_1_1_1_15,
  input      [7:0]    push_payload_1_1_2_0,
  input      [7:0]    push_payload_1_1_2_1,
  input      [7:0]    push_payload_1_1_2_2,
  input      [7:0]    push_payload_1_1_2_3,
  input      [7:0]    push_payload_1_1_2_4,
  input      [7:0]    push_payload_1_1_2_5,
  input      [7:0]    push_payload_1_1_2_6,
  input      [7:0]    push_payload_1_1_2_7,
  input      [7:0]    push_payload_1_1_2_8,
  input      [7:0]    push_payload_1_1_2_9,
  input      [7:0]    push_payload_1_1_2_10,
  input      [7:0]    push_payload_1_1_2_11,
  input      [7:0]    push_payload_1_1_2_12,
  input      [7:0]    push_payload_1_1_2_13,
  input      [7:0]    push_payload_1_1_2_14,
  input      [7:0]    push_payload_1_1_2_15,
  input      [7:0]    push_payload_1_2_0_0,
  input      [7:0]    push_payload_1_2_0_1,
  input      [7:0]    push_payload_1_2_0_2,
  input      [7:0]    push_payload_1_2_0_3,
  input      [7:0]    push_payload_1_2_0_4,
  input      [7:0]    push_payload_1_2_0_5,
  input      [7:0]    push_payload_1_2_0_6,
  input      [7:0]    push_payload_1_2_0_7,
  input      [7:0]    push_payload_1_2_0_8,
  input      [7:0]    push_payload_1_2_0_9,
  input      [7:0]    push_payload_1_2_0_10,
  input      [7:0]    push_payload_1_2_0_11,
  input      [7:0]    push_payload_1_2_0_12,
  input      [7:0]    push_payload_1_2_0_13,
  input      [7:0]    push_payload_1_2_0_14,
  input      [7:0]    push_payload_1_2_0_15,
  input      [7:0]    push_payload_1_2_1_0,
  input      [7:0]    push_payload_1_2_1_1,
  input      [7:0]    push_payload_1_2_1_2,
  input      [7:0]    push_payload_1_2_1_3,
  input      [7:0]    push_payload_1_2_1_4,
  input      [7:0]    push_payload_1_2_1_5,
  input      [7:0]    push_payload_1_2_1_6,
  input      [7:0]    push_payload_1_2_1_7,
  input      [7:0]    push_payload_1_2_1_8,
  input      [7:0]    push_payload_1_2_1_9,
  input      [7:0]    push_payload_1_2_1_10,
  input      [7:0]    push_payload_1_2_1_11,
  input      [7:0]    push_payload_1_2_1_12,
  input      [7:0]    push_payload_1_2_1_13,
  input      [7:0]    push_payload_1_2_1_14,
  input      [7:0]    push_payload_1_2_1_15,
  input      [7:0]    push_payload_1_2_2_0,
  input      [7:0]    push_payload_1_2_2_1,
  input      [7:0]    push_payload_1_2_2_2,
  input      [7:0]    push_payload_1_2_2_3,
  input      [7:0]    push_payload_1_2_2_4,
  input      [7:0]    push_payload_1_2_2_5,
  input      [7:0]    push_payload_1_2_2_6,
  input      [7:0]    push_payload_1_2_2_7,
  input      [7:0]    push_payload_1_2_2_8,
  input      [7:0]    push_payload_1_2_2_9,
  input      [7:0]    push_payload_1_2_2_10,
  input      [7:0]    push_payload_1_2_2_11,
  input      [7:0]    push_payload_1_2_2_12,
  input      [7:0]    push_payload_1_2_2_13,
  input      [7:0]    push_payload_1_2_2_14,
  input      [7:0]    push_payload_1_2_2_15,
  output              pop_valid,
  input               pop_ready,
  output     [7:0]    pop_payload_0_0_0_0,
  output     [7:0]    pop_payload_0_0_0_1,
  output     [7:0]    pop_payload_0_0_0_2,
  output     [7:0]    pop_payload_0_0_0_3,
  output     [7:0]    pop_payload_0_0_0_4,
  output     [7:0]    pop_payload_0_0_0_5,
  output     [7:0]    pop_payload_0_0_0_6,
  output     [7:0]    pop_payload_0_0_0_7,
  output     [7:0]    pop_payload_0_0_0_8,
  output     [7:0]    pop_payload_0_0_0_9,
  output     [7:0]    pop_payload_0_0_0_10,
  output     [7:0]    pop_payload_0_0_0_11,
  output     [7:0]    pop_payload_0_0_0_12,
  output     [7:0]    pop_payload_0_0_0_13,
  output     [7:0]    pop_payload_0_0_0_14,
  output     [7:0]    pop_payload_0_0_0_15,
  output     [7:0]    pop_payload_0_0_1_0,
  output     [7:0]    pop_payload_0_0_1_1,
  output     [7:0]    pop_payload_0_0_1_2,
  output     [7:0]    pop_payload_0_0_1_3,
  output     [7:0]    pop_payload_0_0_1_4,
  output     [7:0]    pop_payload_0_0_1_5,
  output     [7:0]    pop_payload_0_0_1_6,
  output     [7:0]    pop_payload_0_0_1_7,
  output     [7:0]    pop_payload_0_0_1_8,
  output     [7:0]    pop_payload_0_0_1_9,
  output     [7:0]    pop_payload_0_0_1_10,
  output     [7:0]    pop_payload_0_0_1_11,
  output     [7:0]    pop_payload_0_0_1_12,
  output     [7:0]    pop_payload_0_0_1_13,
  output     [7:0]    pop_payload_0_0_1_14,
  output     [7:0]    pop_payload_0_0_1_15,
  output     [7:0]    pop_payload_0_0_2_0,
  output     [7:0]    pop_payload_0_0_2_1,
  output     [7:0]    pop_payload_0_0_2_2,
  output     [7:0]    pop_payload_0_0_2_3,
  output     [7:0]    pop_payload_0_0_2_4,
  output     [7:0]    pop_payload_0_0_2_5,
  output     [7:0]    pop_payload_0_0_2_6,
  output     [7:0]    pop_payload_0_0_2_7,
  output     [7:0]    pop_payload_0_0_2_8,
  output     [7:0]    pop_payload_0_0_2_9,
  output     [7:0]    pop_payload_0_0_2_10,
  output     [7:0]    pop_payload_0_0_2_11,
  output     [7:0]    pop_payload_0_0_2_12,
  output     [7:0]    pop_payload_0_0_2_13,
  output     [7:0]    pop_payload_0_0_2_14,
  output     [7:0]    pop_payload_0_0_2_15,
  output     [7:0]    pop_payload_0_1_0_0,
  output     [7:0]    pop_payload_0_1_0_1,
  output     [7:0]    pop_payload_0_1_0_2,
  output     [7:0]    pop_payload_0_1_0_3,
  output     [7:0]    pop_payload_0_1_0_4,
  output     [7:0]    pop_payload_0_1_0_5,
  output     [7:0]    pop_payload_0_1_0_6,
  output     [7:0]    pop_payload_0_1_0_7,
  output     [7:0]    pop_payload_0_1_0_8,
  output     [7:0]    pop_payload_0_1_0_9,
  output     [7:0]    pop_payload_0_1_0_10,
  output     [7:0]    pop_payload_0_1_0_11,
  output     [7:0]    pop_payload_0_1_0_12,
  output     [7:0]    pop_payload_0_1_0_13,
  output     [7:0]    pop_payload_0_1_0_14,
  output     [7:0]    pop_payload_0_1_0_15,
  output     [7:0]    pop_payload_0_1_1_0,
  output     [7:0]    pop_payload_0_1_1_1,
  output     [7:0]    pop_payload_0_1_1_2,
  output     [7:0]    pop_payload_0_1_1_3,
  output     [7:0]    pop_payload_0_1_1_4,
  output     [7:0]    pop_payload_0_1_1_5,
  output     [7:0]    pop_payload_0_1_1_6,
  output     [7:0]    pop_payload_0_1_1_7,
  output     [7:0]    pop_payload_0_1_1_8,
  output     [7:0]    pop_payload_0_1_1_9,
  output     [7:0]    pop_payload_0_1_1_10,
  output     [7:0]    pop_payload_0_1_1_11,
  output     [7:0]    pop_payload_0_1_1_12,
  output     [7:0]    pop_payload_0_1_1_13,
  output     [7:0]    pop_payload_0_1_1_14,
  output     [7:0]    pop_payload_0_1_1_15,
  output     [7:0]    pop_payload_0_1_2_0,
  output     [7:0]    pop_payload_0_1_2_1,
  output     [7:0]    pop_payload_0_1_2_2,
  output     [7:0]    pop_payload_0_1_2_3,
  output     [7:0]    pop_payload_0_1_2_4,
  output     [7:0]    pop_payload_0_1_2_5,
  output     [7:0]    pop_payload_0_1_2_6,
  output     [7:0]    pop_payload_0_1_2_7,
  output     [7:0]    pop_payload_0_1_2_8,
  output     [7:0]    pop_payload_0_1_2_9,
  output     [7:0]    pop_payload_0_1_2_10,
  output     [7:0]    pop_payload_0_1_2_11,
  output     [7:0]    pop_payload_0_1_2_12,
  output     [7:0]    pop_payload_0_1_2_13,
  output     [7:0]    pop_payload_0_1_2_14,
  output     [7:0]    pop_payload_0_1_2_15,
  output     [7:0]    pop_payload_0_2_0_0,
  output     [7:0]    pop_payload_0_2_0_1,
  output     [7:0]    pop_payload_0_2_0_2,
  output     [7:0]    pop_payload_0_2_0_3,
  output     [7:0]    pop_payload_0_2_0_4,
  output     [7:0]    pop_payload_0_2_0_5,
  output     [7:0]    pop_payload_0_2_0_6,
  output     [7:0]    pop_payload_0_2_0_7,
  output     [7:0]    pop_payload_0_2_0_8,
  output     [7:0]    pop_payload_0_2_0_9,
  output     [7:0]    pop_payload_0_2_0_10,
  output     [7:0]    pop_payload_0_2_0_11,
  output     [7:0]    pop_payload_0_2_0_12,
  output     [7:0]    pop_payload_0_2_0_13,
  output     [7:0]    pop_payload_0_2_0_14,
  output     [7:0]    pop_payload_0_2_0_15,
  output     [7:0]    pop_payload_0_2_1_0,
  output     [7:0]    pop_payload_0_2_1_1,
  output     [7:0]    pop_payload_0_2_1_2,
  output     [7:0]    pop_payload_0_2_1_3,
  output     [7:0]    pop_payload_0_2_1_4,
  output     [7:0]    pop_payload_0_2_1_5,
  output     [7:0]    pop_payload_0_2_1_6,
  output     [7:0]    pop_payload_0_2_1_7,
  output     [7:0]    pop_payload_0_2_1_8,
  output     [7:0]    pop_payload_0_2_1_9,
  output     [7:0]    pop_payload_0_2_1_10,
  output     [7:0]    pop_payload_0_2_1_11,
  output     [7:0]    pop_payload_0_2_1_12,
  output     [7:0]    pop_payload_0_2_1_13,
  output     [7:0]    pop_payload_0_2_1_14,
  output     [7:0]    pop_payload_0_2_1_15,
  output     [7:0]    pop_payload_0_2_2_0,
  output     [7:0]    pop_payload_0_2_2_1,
  output     [7:0]    pop_payload_0_2_2_2,
  output     [7:0]    pop_payload_0_2_2_3,
  output     [7:0]    pop_payload_0_2_2_4,
  output     [7:0]    pop_payload_0_2_2_5,
  output     [7:0]    pop_payload_0_2_2_6,
  output     [7:0]    pop_payload_0_2_2_7,
  output     [7:0]    pop_payload_0_2_2_8,
  output     [7:0]    pop_payload_0_2_2_9,
  output     [7:0]    pop_payload_0_2_2_10,
  output     [7:0]    pop_payload_0_2_2_11,
  output     [7:0]    pop_payload_0_2_2_12,
  output     [7:0]    pop_payload_0_2_2_13,
  output     [7:0]    pop_payload_0_2_2_14,
  output     [7:0]    pop_payload_0_2_2_15,
  output     [7:0]    pop_payload_1_0_0_0,
  output     [7:0]    pop_payload_1_0_0_1,
  output     [7:0]    pop_payload_1_0_0_2,
  output     [7:0]    pop_payload_1_0_0_3,
  output     [7:0]    pop_payload_1_0_0_4,
  output     [7:0]    pop_payload_1_0_0_5,
  output     [7:0]    pop_payload_1_0_0_6,
  output     [7:0]    pop_payload_1_0_0_7,
  output     [7:0]    pop_payload_1_0_0_8,
  output     [7:0]    pop_payload_1_0_0_9,
  output     [7:0]    pop_payload_1_0_0_10,
  output     [7:0]    pop_payload_1_0_0_11,
  output     [7:0]    pop_payload_1_0_0_12,
  output     [7:0]    pop_payload_1_0_0_13,
  output     [7:0]    pop_payload_1_0_0_14,
  output     [7:0]    pop_payload_1_0_0_15,
  output     [7:0]    pop_payload_1_0_1_0,
  output     [7:0]    pop_payload_1_0_1_1,
  output     [7:0]    pop_payload_1_0_1_2,
  output     [7:0]    pop_payload_1_0_1_3,
  output     [7:0]    pop_payload_1_0_1_4,
  output     [7:0]    pop_payload_1_0_1_5,
  output     [7:0]    pop_payload_1_0_1_6,
  output     [7:0]    pop_payload_1_0_1_7,
  output     [7:0]    pop_payload_1_0_1_8,
  output     [7:0]    pop_payload_1_0_1_9,
  output     [7:0]    pop_payload_1_0_1_10,
  output     [7:0]    pop_payload_1_0_1_11,
  output     [7:0]    pop_payload_1_0_1_12,
  output     [7:0]    pop_payload_1_0_1_13,
  output     [7:0]    pop_payload_1_0_1_14,
  output     [7:0]    pop_payload_1_0_1_15,
  output     [7:0]    pop_payload_1_0_2_0,
  output     [7:0]    pop_payload_1_0_2_1,
  output     [7:0]    pop_payload_1_0_2_2,
  output     [7:0]    pop_payload_1_0_2_3,
  output     [7:0]    pop_payload_1_0_2_4,
  output     [7:0]    pop_payload_1_0_2_5,
  output     [7:0]    pop_payload_1_0_2_6,
  output     [7:0]    pop_payload_1_0_2_7,
  output     [7:0]    pop_payload_1_0_2_8,
  output     [7:0]    pop_payload_1_0_2_9,
  output     [7:0]    pop_payload_1_0_2_10,
  output     [7:0]    pop_payload_1_0_2_11,
  output     [7:0]    pop_payload_1_0_2_12,
  output     [7:0]    pop_payload_1_0_2_13,
  output     [7:0]    pop_payload_1_0_2_14,
  output     [7:0]    pop_payload_1_0_2_15,
  output     [7:0]    pop_payload_1_1_0_0,
  output     [7:0]    pop_payload_1_1_0_1,
  output     [7:0]    pop_payload_1_1_0_2,
  output     [7:0]    pop_payload_1_1_0_3,
  output     [7:0]    pop_payload_1_1_0_4,
  output     [7:0]    pop_payload_1_1_0_5,
  output     [7:0]    pop_payload_1_1_0_6,
  output     [7:0]    pop_payload_1_1_0_7,
  output     [7:0]    pop_payload_1_1_0_8,
  output     [7:0]    pop_payload_1_1_0_9,
  output     [7:0]    pop_payload_1_1_0_10,
  output     [7:0]    pop_payload_1_1_0_11,
  output     [7:0]    pop_payload_1_1_0_12,
  output     [7:0]    pop_payload_1_1_0_13,
  output     [7:0]    pop_payload_1_1_0_14,
  output     [7:0]    pop_payload_1_1_0_15,
  output     [7:0]    pop_payload_1_1_1_0,
  output     [7:0]    pop_payload_1_1_1_1,
  output     [7:0]    pop_payload_1_1_1_2,
  output     [7:0]    pop_payload_1_1_1_3,
  output     [7:0]    pop_payload_1_1_1_4,
  output     [7:0]    pop_payload_1_1_1_5,
  output     [7:0]    pop_payload_1_1_1_6,
  output     [7:0]    pop_payload_1_1_1_7,
  output     [7:0]    pop_payload_1_1_1_8,
  output     [7:0]    pop_payload_1_1_1_9,
  output     [7:0]    pop_payload_1_1_1_10,
  output     [7:0]    pop_payload_1_1_1_11,
  output     [7:0]    pop_payload_1_1_1_12,
  output     [7:0]    pop_payload_1_1_1_13,
  output     [7:0]    pop_payload_1_1_1_14,
  output     [7:0]    pop_payload_1_1_1_15,
  output     [7:0]    pop_payload_1_1_2_0,
  output     [7:0]    pop_payload_1_1_2_1,
  output     [7:0]    pop_payload_1_1_2_2,
  output     [7:0]    pop_payload_1_1_2_3,
  output     [7:0]    pop_payload_1_1_2_4,
  output     [7:0]    pop_payload_1_1_2_5,
  output     [7:0]    pop_payload_1_1_2_6,
  output     [7:0]    pop_payload_1_1_2_7,
  output     [7:0]    pop_payload_1_1_2_8,
  output     [7:0]    pop_payload_1_1_2_9,
  output     [7:0]    pop_payload_1_1_2_10,
  output     [7:0]    pop_payload_1_1_2_11,
  output     [7:0]    pop_payload_1_1_2_12,
  output     [7:0]    pop_payload_1_1_2_13,
  output     [7:0]    pop_payload_1_1_2_14,
  output     [7:0]    pop_payload_1_1_2_15,
  output     [7:0]    pop_payload_1_2_0_0,
  output     [7:0]    pop_payload_1_2_0_1,
  output     [7:0]    pop_payload_1_2_0_2,
  output     [7:0]    pop_payload_1_2_0_3,
  output     [7:0]    pop_payload_1_2_0_4,
  output     [7:0]    pop_payload_1_2_0_5,
  output     [7:0]    pop_payload_1_2_0_6,
  output     [7:0]    pop_payload_1_2_0_7,
  output     [7:0]    pop_payload_1_2_0_8,
  output     [7:0]    pop_payload_1_2_0_9,
  output     [7:0]    pop_payload_1_2_0_10,
  output     [7:0]    pop_payload_1_2_0_11,
  output     [7:0]    pop_payload_1_2_0_12,
  output     [7:0]    pop_payload_1_2_0_13,
  output     [7:0]    pop_payload_1_2_0_14,
  output     [7:0]    pop_payload_1_2_0_15,
  output     [7:0]    pop_payload_1_2_1_0,
  output     [7:0]    pop_payload_1_2_1_1,
  output     [7:0]    pop_payload_1_2_1_2,
  output     [7:0]    pop_payload_1_2_1_3,
  output     [7:0]    pop_payload_1_2_1_4,
  output     [7:0]    pop_payload_1_2_1_5,
  output     [7:0]    pop_payload_1_2_1_6,
  output     [7:0]    pop_payload_1_2_1_7,
  output     [7:0]    pop_payload_1_2_1_8,
  output     [7:0]    pop_payload_1_2_1_9,
  output     [7:0]    pop_payload_1_2_1_10,
  output     [7:0]    pop_payload_1_2_1_11,
  output     [7:0]    pop_payload_1_2_1_12,
  output     [7:0]    pop_payload_1_2_1_13,
  output     [7:0]    pop_payload_1_2_1_14,
  output     [7:0]    pop_payload_1_2_1_15,
  output     [7:0]    pop_payload_1_2_2_0,
  output     [7:0]    pop_payload_1_2_2_1,
  output     [7:0]    pop_payload_1_2_2_2,
  output     [7:0]    pop_payload_1_2_2_3,
  output     [7:0]    pop_payload_1_2_2_4,
  output     [7:0]    pop_payload_1_2_2_5,
  output     [7:0]    pop_payload_1_2_2_6,
  output     [7:0]    pop_payload_1_2_2_7,
  output     [7:0]    pop_payload_1_2_2_8,
  output     [7:0]    pop_payload_1_2_2_9,
  output     [7:0]    pop_payload_1_2_2_10,
  output     [7:0]    pop_payload_1_2_2_11,
  output     [7:0]    pop_payload_1_2_2_12,
  output     [7:0]    pop_payload_1_2_2_13,
  output     [7:0]    pop_payload_1_2_2_14,
  output     [7:0]    pop_payload_1_2_2_15,
  input               flush,
  input               clk,
  input               reset
);

  reg        [2303:0] tmp_ram_port0;
  wire       [4:0]    tmp_pushPtr_valueNext;
  wire       [0:0]    tmp_pushPtr_valueNext_1;
  wire       [4:0]    tmp_popPtr_valueNext;
  wire       [0:0]    tmp_popPtr_valueNext_1;
  wire       [2303:0] tmp_ram_port;
  reg                 tmp_1;
  wire                popEvent_valid;
  reg                 popEvent_ready;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [4:0]    pushPtr_valueNext;
  reg        [4:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [4:0]    popPtr_valueNext;
  reg        [4:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                pushing;
  wire                popping;
  wire                empty;
  wire                full;
  reg                 tmp_popEvent_valid;
  reg                 rValid;
  wire       [7:0]    rData_0_0_0_0;
  wire       [7:0]    rData_0_0_0_1;
  wire       [7:0]    rData_0_0_0_2;
  wire       [7:0]    rData_0_0_0_3;
  wire       [7:0]    rData_0_0_0_4;
  wire       [7:0]    rData_0_0_0_5;
  wire       [7:0]    rData_0_0_0_6;
  wire       [7:0]    rData_0_0_0_7;
  wire       [7:0]    rData_0_0_0_8;
  wire       [7:0]    rData_0_0_0_9;
  wire       [7:0]    rData_0_0_0_10;
  wire       [7:0]    rData_0_0_0_11;
  wire       [7:0]    rData_0_0_0_12;
  wire       [7:0]    rData_0_0_0_13;
  wire       [7:0]    rData_0_0_0_14;
  wire       [7:0]    rData_0_0_0_15;
  wire       [7:0]    rData_0_0_1_0;
  wire       [7:0]    rData_0_0_1_1;
  wire       [7:0]    rData_0_0_1_2;
  wire       [7:0]    rData_0_0_1_3;
  wire       [7:0]    rData_0_0_1_4;
  wire       [7:0]    rData_0_0_1_5;
  wire       [7:0]    rData_0_0_1_6;
  wire       [7:0]    rData_0_0_1_7;
  wire       [7:0]    rData_0_0_1_8;
  wire       [7:0]    rData_0_0_1_9;
  wire       [7:0]    rData_0_0_1_10;
  wire       [7:0]    rData_0_0_1_11;
  wire       [7:0]    rData_0_0_1_12;
  wire       [7:0]    rData_0_0_1_13;
  wire       [7:0]    rData_0_0_1_14;
  wire       [7:0]    rData_0_0_1_15;
  wire       [7:0]    rData_0_0_2_0;
  wire       [7:0]    rData_0_0_2_1;
  wire       [7:0]    rData_0_0_2_2;
  wire       [7:0]    rData_0_0_2_3;
  wire       [7:0]    rData_0_0_2_4;
  wire       [7:0]    rData_0_0_2_5;
  wire       [7:0]    rData_0_0_2_6;
  wire       [7:0]    rData_0_0_2_7;
  wire       [7:0]    rData_0_0_2_8;
  wire       [7:0]    rData_0_0_2_9;
  wire       [7:0]    rData_0_0_2_10;
  wire       [7:0]    rData_0_0_2_11;
  wire       [7:0]    rData_0_0_2_12;
  wire       [7:0]    rData_0_0_2_13;
  wire       [7:0]    rData_0_0_2_14;
  wire       [7:0]    rData_0_0_2_15;
  wire       [7:0]    rData_0_1_0_0;
  wire       [7:0]    rData_0_1_0_1;
  wire       [7:0]    rData_0_1_0_2;
  wire       [7:0]    rData_0_1_0_3;
  wire       [7:0]    rData_0_1_0_4;
  wire       [7:0]    rData_0_1_0_5;
  wire       [7:0]    rData_0_1_0_6;
  wire       [7:0]    rData_0_1_0_7;
  wire       [7:0]    rData_0_1_0_8;
  wire       [7:0]    rData_0_1_0_9;
  wire       [7:0]    rData_0_1_0_10;
  wire       [7:0]    rData_0_1_0_11;
  wire       [7:0]    rData_0_1_0_12;
  wire       [7:0]    rData_0_1_0_13;
  wire       [7:0]    rData_0_1_0_14;
  wire       [7:0]    rData_0_1_0_15;
  wire       [7:0]    rData_0_1_1_0;
  wire       [7:0]    rData_0_1_1_1;
  wire       [7:0]    rData_0_1_1_2;
  wire       [7:0]    rData_0_1_1_3;
  wire       [7:0]    rData_0_1_1_4;
  wire       [7:0]    rData_0_1_1_5;
  wire       [7:0]    rData_0_1_1_6;
  wire       [7:0]    rData_0_1_1_7;
  wire       [7:0]    rData_0_1_1_8;
  wire       [7:0]    rData_0_1_1_9;
  wire       [7:0]    rData_0_1_1_10;
  wire       [7:0]    rData_0_1_1_11;
  wire       [7:0]    rData_0_1_1_12;
  wire       [7:0]    rData_0_1_1_13;
  wire       [7:0]    rData_0_1_1_14;
  wire       [7:0]    rData_0_1_1_15;
  wire       [7:0]    rData_0_1_2_0;
  wire       [7:0]    rData_0_1_2_1;
  wire       [7:0]    rData_0_1_2_2;
  wire       [7:0]    rData_0_1_2_3;
  wire       [7:0]    rData_0_1_2_4;
  wire       [7:0]    rData_0_1_2_5;
  wire       [7:0]    rData_0_1_2_6;
  wire       [7:0]    rData_0_1_2_7;
  wire       [7:0]    rData_0_1_2_8;
  wire       [7:0]    rData_0_1_2_9;
  wire       [7:0]    rData_0_1_2_10;
  wire       [7:0]    rData_0_1_2_11;
  wire       [7:0]    rData_0_1_2_12;
  wire       [7:0]    rData_0_1_2_13;
  wire       [7:0]    rData_0_1_2_14;
  wire       [7:0]    rData_0_1_2_15;
  wire       [7:0]    rData_0_2_0_0;
  wire       [7:0]    rData_0_2_0_1;
  wire       [7:0]    rData_0_2_0_2;
  wire       [7:0]    rData_0_2_0_3;
  wire       [7:0]    rData_0_2_0_4;
  wire       [7:0]    rData_0_2_0_5;
  wire       [7:0]    rData_0_2_0_6;
  wire       [7:0]    rData_0_2_0_7;
  wire       [7:0]    rData_0_2_0_8;
  wire       [7:0]    rData_0_2_0_9;
  wire       [7:0]    rData_0_2_0_10;
  wire       [7:0]    rData_0_2_0_11;
  wire       [7:0]    rData_0_2_0_12;
  wire       [7:0]    rData_0_2_0_13;
  wire       [7:0]    rData_0_2_0_14;
  wire       [7:0]    rData_0_2_0_15;
  wire       [7:0]    rData_0_2_1_0;
  wire       [7:0]    rData_0_2_1_1;
  wire       [7:0]    rData_0_2_1_2;
  wire       [7:0]    rData_0_2_1_3;
  wire       [7:0]    rData_0_2_1_4;
  wire       [7:0]    rData_0_2_1_5;
  wire       [7:0]    rData_0_2_1_6;
  wire       [7:0]    rData_0_2_1_7;
  wire       [7:0]    rData_0_2_1_8;
  wire       [7:0]    rData_0_2_1_9;
  wire       [7:0]    rData_0_2_1_10;
  wire       [7:0]    rData_0_2_1_11;
  wire       [7:0]    rData_0_2_1_12;
  wire       [7:0]    rData_0_2_1_13;
  wire       [7:0]    rData_0_2_1_14;
  wire       [7:0]    rData_0_2_1_15;
  wire       [7:0]    rData_0_2_2_0;
  wire       [7:0]    rData_0_2_2_1;
  wire       [7:0]    rData_0_2_2_2;
  wire       [7:0]    rData_0_2_2_3;
  wire       [7:0]    rData_0_2_2_4;
  wire       [7:0]    rData_0_2_2_5;
  wire       [7:0]    rData_0_2_2_6;
  wire       [7:0]    rData_0_2_2_7;
  wire       [7:0]    rData_0_2_2_8;
  wire       [7:0]    rData_0_2_2_9;
  wire       [7:0]    rData_0_2_2_10;
  wire       [7:0]    rData_0_2_2_11;
  wire       [7:0]    rData_0_2_2_12;
  wire       [7:0]    rData_0_2_2_13;
  wire       [7:0]    rData_0_2_2_14;
  wire       [7:0]    rData_0_2_2_15;
  wire       [7:0]    rData_1_0_0_0;
  wire       [7:0]    rData_1_0_0_1;
  wire       [7:0]    rData_1_0_0_2;
  wire       [7:0]    rData_1_0_0_3;
  wire       [7:0]    rData_1_0_0_4;
  wire       [7:0]    rData_1_0_0_5;
  wire       [7:0]    rData_1_0_0_6;
  wire       [7:0]    rData_1_0_0_7;
  wire       [7:0]    rData_1_0_0_8;
  wire       [7:0]    rData_1_0_0_9;
  wire       [7:0]    rData_1_0_0_10;
  wire       [7:0]    rData_1_0_0_11;
  wire       [7:0]    rData_1_0_0_12;
  wire       [7:0]    rData_1_0_0_13;
  wire       [7:0]    rData_1_0_0_14;
  wire       [7:0]    rData_1_0_0_15;
  wire       [7:0]    rData_1_0_1_0;
  wire       [7:0]    rData_1_0_1_1;
  wire       [7:0]    rData_1_0_1_2;
  wire       [7:0]    rData_1_0_1_3;
  wire       [7:0]    rData_1_0_1_4;
  wire       [7:0]    rData_1_0_1_5;
  wire       [7:0]    rData_1_0_1_6;
  wire       [7:0]    rData_1_0_1_7;
  wire       [7:0]    rData_1_0_1_8;
  wire       [7:0]    rData_1_0_1_9;
  wire       [7:0]    rData_1_0_1_10;
  wire       [7:0]    rData_1_0_1_11;
  wire       [7:0]    rData_1_0_1_12;
  wire       [7:0]    rData_1_0_1_13;
  wire       [7:0]    rData_1_0_1_14;
  wire       [7:0]    rData_1_0_1_15;
  wire       [7:0]    rData_1_0_2_0;
  wire       [7:0]    rData_1_0_2_1;
  wire       [7:0]    rData_1_0_2_2;
  wire       [7:0]    rData_1_0_2_3;
  wire       [7:0]    rData_1_0_2_4;
  wire       [7:0]    rData_1_0_2_5;
  wire       [7:0]    rData_1_0_2_6;
  wire       [7:0]    rData_1_0_2_7;
  wire       [7:0]    rData_1_0_2_8;
  wire       [7:0]    rData_1_0_2_9;
  wire       [7:0]    rData_1_0_2_10;
  wire       [7:0]    rData_1_0_2_11;
  wire       [7:0]    rData_1_0_2_12;
  wire       [7:0]    rData_1_0_2_13;
  wire       [7:0]    rData_1_0_2_14;
  wire       [7:0]    rData_1_0_2_15;
  wire       [7:0]    rData_1_1_0_0;
  wire       [7:0]    rData_1_1_0_1;
  wire       [7:0]    rData_1_1_0_2;
  wire       [7:0]    rData_1_1_0_3;
  wire       [7:0]    rData_1_1_0_4;
  wire       [7:0]    rData_1_1_0_5;
  wire       [7:0]    rData_1_1_0_6;
  wire       [7:0]    rData_1_1_0_7;
  wire       [7:0]    rData_1_1_0_8;
  wire       [7:0]    rData_1_1_0_9;
  wire       [7:0]    rData_1_1_0_10;
  wire       [7:0]    rData_1_1_0_11;
  wire       [7:0]    rData_1_1_0_12;
  wire       [7:0]    rData_1_1_0_13;
  wire       [7:0]    rData_1_1_0_14;
  wire       [7:0]    rData_1_1_0_15;
  wire       [7:0]    rData_1_1_1_0;
  wire       [7:0]    rData_1_1_1_1;
  wire       [7:0]    rData_1_1_1_2;
  wire       [7:0]    rData_1_1_1_3;
  wire       [7:0]    rData_1_1_1_4;
  wire       [7:0]    rData_1_1_1_5;
  wire       [7:0]    rData_1_1_1_6;
  wire       [7:0]    rData_1_1_1_7;
  wire       [7:0]    rData_1_1_1_8;
  wire       [7:0]    rData_1_1_1_9;
  wire       [7:0]    rData_1_1_1_10;
  wire       [7:0]    rData_1_1_1_11;
  wire       [7:0]    rData_1_1_1_12;
  wire       [7:0]    rData_1_1_1_13;
  wire       [7:0]    rData_1_1_1_14;
  wire       [7:0]    rData_1_1_1_15;
  wire       [7:0]    rData_1_1_2_0;
  wire       [7:0]    rData_1_1_2_1;
  wire       [7:0]    rData_1_1_2_2;
  wire       [7:0]    rData_1_1_2_3;
  wire       [7:0]    rData_1_1_2_4;
  wire       [7:0]    rData_1_1_2_5;
  wire       [7:0]    rData_1_1_2_6;
  wire       [7:0]    rData_1_1_2_7;
  wire       [7:0]    rData_1_1_2_8;
  wire       [7:0]    rData_1_1_2_9;
  wire       [7:0]    rData_1_1_2_10;
  wire       [7:0]    rData_1_1_2_11;
  wire       [7:0]    rData_1_1_2_12;
  wire       [7:0]    rData_1_1_2_13;
  wire       [7:0]    rData_1_1_2_14;
  wire       [7:0]    rData_1_1_2_15;
  wire       [7:0]    rData_1_2_0_0;
  wire       [7:0]    rData_1_2_0_1;
  wire       [7:0]    rData_1_2_0_2;
  wire       [7:0]    rData_1_2_0_3;
  wire       [7:0]    rData_1_2_0_4;
  wire       [7:0]    rData_1_2_0_5;
  wire       [7:0]    rData_1_2_0_6;
  wire       [7:0]    rData_1_2_0_7;
  wire       [7:0]    rData_1_2_0_8;
  wire       [7:0]    rData_1_2_0_9;
  wire       [7:0]    rData_1_2_0_10;
  wire       [7:0]    rData_1_2_0_11;
  wire       [7:0]    rData_1_2_0_12;
  wire       [7:0]    rData_1_2_0_13;
  wire       [7:0]    rData_1_2_0_14;
  wire       [7:0]    rData_1_2_0_15;
  wire       [7:0]    rData_1_2_1_0;
  wire       [7:0]    rData_1_2_1_1;
  wire       [7:0]    rData_1_2_1_2;
  wire       [7:0]    rData_1_2_1_3;
  wire       [7:0]    rData_1_2_1_4;
  wire       [7:0]    rData_1_2_1_5;
  wire       [7:0]    rData_1_2_1_6;
  wire       [7:0]    rData_1_2_1_7;
  wire       [7:0]    rData_1_2_1_8;
  wire       [7:0]    rData_1_2_1_9;
  wire       [7:0]    rData_1_2_1_10;
  wire       [7:0]    rData_1_2_1_11;
  wire       [7:0]    rData_1_2_1_12;
  wire       [7:0]    rData_1_2_1_13;
  wire       [7:0]    rData_1_2_1_14;
  wire       [7:0]    rData_1_2_1_15;
  wire       [7:0]    rData_1_2_2_0;
  wire       [7:0]    rData_1_2_2_1;
  wire       [7:0]    rData_1_2_2_2;
  wire       [7:0]    rData_1_2_2_3;
  wire       [7:0]    rData_1_2_2_4;
  wire       [7:0]    rData_1_2_2_5;
  wire       [7:0]    rData_1_2_2_6;
  wire       [7:0]    rData_1_2_2_7;
  wire       [7:0]    rData_1_2_2_8;
  wire       [7:0]    rData_1_2_2_9;
  wire       [7:0]    rData_1_2_2_10;
  wire       [7:0]    rData_1_2_2_11;
  wire       [7:0]    rData_1_2_2_12;
  wire       [7:0]    rData_1_2_2_13;
  wire       [7:0]    rData_1_2_2_14;
  wire       [7:0]    rData_1_2_2_15;
  wire       [2303:0] tmp_rData_0_0_0_0;
  wire       [1151:0] tmp_rData_0_0_0_0_1;
  wire       [383:0]  tmp_rData_0_0_0_0_2;
  wire       [127:0]  tmp_rData_0_0_0_0_3;
  wire       [127:0]  tmp_rData_0_0_1_0;
  wire       [127:0]  tmp_rData_0_0_2_0;
  wire       [383:0]  tmp_rData_0_1_0_0;
  wire       [127:0]  tmp_rData_0_1_0_0_1;
  wire       [127:0]  tmp_rData_0_1_1_0;
  wire       [127:0]  tmp_rData_0_1_2_0;
  wire       [383:0]  tmp_rData_0_2_0_0;
  wire       [127:0]  tmp_rData_0_2_0_0_1;
  wire       [127:0]  tmp_rData_0_2_1_0;
  wire       [127:0]  tmp_rData_0_2_2_0;
  wire       [1151:0] tmp_rData_1_0_0_0;
  wire       [383:0]  tmp_rData_1_0_0_0_1;
  wire       [127:0]  tmp_rData_1_0_0_0_2;
  wire       [127:0]  tmp_rData_1_0_1_0;
  wire       [127:0]  tmp_rData_1_0_2_0;
  wire       [383:0]  tmp_rData_1_1_0_0;
  wire       [127:0]  tmp_rData_1_1_0_0_1;
  wire       [127:0]  tmp_rData_1_1_1_0;
  wire       [127:0]  tmp_rData_1_1_2_0;
  wire       [383:0]  tmp_rData_1_2_0_0;
  wire       [127:0]  tmp_rData_1_2_0_0_1;
  wire       [127:0]  tmp_rData_1_2_1_0;
  wire       [127:0]  tmp_rData_1_2_2_0;
  wire                when_StreamFifoHighPerf_l38;
  wire                when_StreamFifoHighPerf_l42;
  (* ram_style = "distributed" *) reg [2303:0] ram [0:31];

  assign tmp_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign tmp_pushPtr_valueNext = {4'd0, tmp_pushPtr_valueNext_1};
  assign tmp_popPtr_valueNext_1 = popPtr_willIncrement;
  assign tmp_popPtr_valueNext = {4'd0, tmp_popPtr_valueNext_1};
  assign tmp_ram_port = {{{{push_payload_1_2_2_15,{push_payload_1_2_2_14,{push_payload_1_2_2_13,{push_payload_1_2_2_12,{push_payload_1_2_2_11,{push_payload_1_2_2_10,{push_payload_1_2_2_9,{push_payload_1_2_2_8,{push_payload_1_2_2_7,{push_payload_1_2_2_6,{push_payload_1_2_2_5,{push_payload_1_2_2_4,{push_payload_1_2_2_3,{push_payload_1_2_2_2,{push_payload_1_2_2_1,push_payload_1_2_2_0}}}}}}}}}}}}}}},{{push_payload_1_2_1_15,{push_payload_1_2_1_14,{push_payload_1_2_1_13,{push_payload_1_2_1_12,{push_payload_1_2_1_11,{push_payload_1_2_1_10,{push_payload_1_2_1_9,{push_payload_1_2_1_8,{push_payload_1_2_1_7,{push_payload_1_2_1_6,{push_payload_1_2_1_5,{push_payload_1_2_1_4,{push_payload_1_2_1_3,{push_payload_1_2_1_2,{push_payload_1_2_1_1,push_payload_1_2_1_0}}}}}}}}}}}}}}},{push_payload_1_2_0_15,{push_payload_1_2_0_14,{push_payload_1_2_0_13,{push_payload_1_2_0_12,{push_payload_1_2_0_11,{push_payload_1_2_0_10,{push_payload_1_2_0_9,{push_payload_1_2_0_8,{push_payload_1_2_0_7,{push_payload_1_2_0_6,{push_payload_1_2_0_5,{push_payload_1_2_0_4,{push_payload_1_2_0_3,{push_payload_1_2_0_2,{push_payload_1_2_0_1,push_payload_1_2_0_0}}}}}}}}}}}}}}}}},{{{push_payload_1_1_2_15,{push_payload_1_1_2_14,{push_payload_1_1_2_13,{push_payload_1_1_2_12,{push_payload_1_1_2_11,{push_payload_1_1_2_10,{push_payload_1_1_2_9,{push_payload_1_1_2_8,{push_payload_1_1_2_7,{push_payload_1_1_2_6,{push_payload_1_1_2_5,{push_payload_1_1_2_4,{push_payload_1_1_2_3,{push_payload_1_1_2_2,{push_payload_1_1_2_1,push_payload_1_1_2_0}}}}}}}}}}}}}}},{{push_payload_1_1_1_15,{push_payload_1_1_1_14,{push_payload_1_1_1_13,{push_payload_1_1_1_12,{push_payload_1_1_1_11,{push_payload_1_1_1_10,{push_payload_1_1_1_9,{push_payload_1_1_1_8,{push_payload_1_1_1_7,{push_payload_1_1_1_6,{push_payload_1_1_1_5,{push_payload_1_1_1_4,{push_payload_1_1_1_3,{push_payload_1_1_1_2,{push_payload_1_1_1_1,push_payload_1_1_1_0}}}}}}}}}}}}}}},{push_payload_1_1_0_15,{push_payload_1_1_0_14,{push_payload_1_1_0_13,{push_payload_1_1_0_12,{push_payload_1_1_0_11,{push_payload_1_1_0_10,{push_payload_1_1_0_9,{push_payload_1_1_0_8,{push_payload_1_1_0_7,{push_payload_1_1_0_6,{push_payload_1_1_0_5,{push_payload_1_1_0_4,{push_payload_1_1_0_3,{push_payload_1_1_0_2,{push_payload_1_1_0_1,push_payload_1_1_0_0}}}}}}}}}}}}}}}}},{{push_payload_1_0_2_15,{push_payload_1_0_2_14,{push_payload_1_0_2_13,{push_payload_1_0_2_12,{push_payload_1_0_2_11,{push_payload_1_0_2_10,{push_payload_1_0_2_9,{push_payload_1_0_2_8,{push_payload_1_0_2_7,{push_payload_1_0_2_6,{push_payload_1_0_2_5,{push_payload_1_0_2_4,{push_payload_1_0_2_3,{push_payload_1_0_2_2,{push_payload_1_0_2_1,push_payload_1_0_2_0}}}}}}}}}}}}}}},{{push_payload_1_0_1_15,{push_payload_1_0_1_14,{push_payload_1_0_1_13,{push_payload_1_0_1_12,{push_payload_1_0_1_11,{push_payload_1_0_1_10,{push_payload_1_0_1_9,{push_payload_1_0_1_8,{push_payload_1_0_1_7,{push_payload_1_0_1_6,{push_payload_1_0_1_5,{push_payload_1_0_1_4,{push_payload_1_0_1_3,{push_payload_1_0_1_2,{push_payload_1_0_1_1,push_payload_1_0_1_0}}}}}}}}}}}}}}},{push_payload_1_0_0_15,{push_payload_1_0_0_14,{push_payload_1_0_0_13,{push_payload_1_0_0_12,{push_payload_1_0_0_11,{push_payload_1_0_0_10,{push_payload_1_0_0_9,{push_payload_1_0_0_8,{push_payload_1_0_0_7,{push_payload_1_0_0_6,{push_payload_1_0_0_5,{push_payload_1_0_0_4,{push_payload_1_0_0_3,{push_payload_1_0_0_2,{push_payload_1_0_0_1,push_payload_1_0_0_0}}}}}}}}}}}}}}}}}}},{{{push_payload_0_2_2_15,{push_payload_0_2_2_14,{push_payload_0_2_2_13,{push_payload_0_2_2_12,{push_payload_0_2_2_11,{push_payload_0_2_2_10,{push_payload_0_2_2_9,{push_payload_0_2_2_8,{push_payload_0_2_2_7,{push_payload_0_2_2_6,{push_payload_0_2_2_5,{push_payload_0_2_2_4,{push_payload_0_2_2_3,{push_payload_0_2_2_2,{push_payload_0_2_2_1,push_payload_0_2_2_0}}}}}}}}}}}}}}},{{push_payload_0_2_1_15,{push_payload_0_2_1_14,{push_payload_0_2_1_13,{push_payload_0_2_1_12,{push_payload_0_2_1_11,{push_payload_0_2_1_10,{push_payload_0_2_1_9,{push_payload_0_2_1_8,{push_payload_0_2_1_7,{push_payload_0_2_1_6,{push_payload_0_2_1_5,{push_payload_0_2_1_4,{push_payload_0_2_1_3,{push_payload_0_2_1_2,{push_payload_0_2_1_1,push_payload_0_2_1_0}}}}}}}}}}}}}}},{push_payload_0_2_0_15,{push_payload_0_2_0_14,{push_payload_0_2_0_13,{push_payload_0_2_0_12,{push_payload_0_2_0_11,{push_payload_0_2_0_10,{push_payload_0_2_0_9,{push_payload_0_2_0_8,{push_payload_0_2_0_7,{push_payload_0_2_0_6,{push_payload_0_2_0_5,{push_payload_0_2_0_4,{push_payload_0_2_0_3,{push_payload_0_2_0_2,{push_payload_0_2_0_1,push_payload_0_2_0_0}}}}}}}}}}}}}}}}},{{{push_payload_0_1_2_15,{push_payload_0_1_2_14,{push_payload_0_1_2_13,{push_payload_0_1_2_12,{push_payload_0_1_2_11,{push_payload_0_1_2_10,{push_payload_0_1_2_9,{push_payload_0_1_2_8,{push_payload_0_1_2_7,{push_payload_0_1_2_6,{push_payload_0_1_2_5,{push_payload_0_1_2_4,{push_payload_0_1_2_3,{push_payload_0_1_2_2,{push_payload_0_1_2_1,push_payload_0_1_2_0}}}}}}}}}}}}}}},{{push_payload_0_1_1_15,{push_payload_0_1_1_14,{push_payload_0_1_1_13,{push_payload_0_1_1_12,{push_payload_0_1_1_11,{push_payload_0_1_1_10,{push_payload_0_1_1_9,{push_payload_0_1_1_8,{push_payload_0_1_1_7,{push_payload_0_1_1_6,{push_payload_0_1_1_5,{push_payload_0_1_1_4,{push_payload_0_1_1_3,{push_payload_0_1_1_2,{push_payload_0_1_1_1,push_payload_0_1_1_0}}}}}}}}}}}}}}},{push_payload_0_1_0_15,{push_payload_0_1_0_14,{push_payload_0_1_0_13,{push_payload_0_1_0_12,{push_payload_0_1_0_11,{push_payload_0_1_0_10,{push_payload_0_1_0_9,{push_payload_0_1_0_8,{push_payload_0_1_0_7,{push_payload_0_1_0_6,{push_payload_0_1_0_5,{push_payload_0_1_0_4,{push_payload_0_1_0_3,{push_payload_0_1_0_2,{push_payload_0_1_0_1,push_payload_0_1_0_0}}}}}}}}}}}}}}}}},{{push_payload_0_0_2_15,{push_payload_0_0_2_14,{push_payload_0_0_2_13,{push_payload_0_0_2_12,{push_payload_0_0_2_11,{push_payload_0_0_2_10,{push_payload_0_0_2_9,{push_payload_0_0_2_8,{push_payload_0_0_2_7,{push_payload_0_0_2_6,{push_payload_0_0_2_5,{push_payload_0_0_2_4,{push_payload_0_0_2_3,{push_payload_0_0_2_2,{push_payload_0_0_2_1,push_payload_0_0_2_0}}}}}}}}}}}}}}},{{push_payload_0_0_1_15,{push_payload_0_0_1_14,{push_payload_0_0_1_13,{push_payload_0_0_1_12,{push_payload_0_0_1_11,{push_payload_0_0_1_10,{push_payload_0_0_1_9,{push_payload_0_0_1_8,{push_payload_0_0_1_7,{push_payload_0_0_1_6,{push_payload_0_0_1_5,{push_payload_0_0_1_4,{push_payload_0_0_1_3,{push_payload_0_0_1_2,{push_payload_0_0_1_1,push_payload_0_0_1_0}}}}}}}}}}}}}}},{push_payload_0_0_0_15,{push_payload_0_0_0_14,{push_payload_0_0_0_13,{push_payload_0_0_0_12,{push_payload_0_0_0_11,{push_payload_0_0_0_10,{push_payload_0_0_0_9,{push_payload_0_0_0_8,{push_payload_0_0_0_7,{push_payload_0_0_0_6,{push_payload_0_0_0_5,{push_payload_0_0_0_4,{push_payload_0_0_0_3,{push_payload_0_0_0_2,{push_payload_0_0_0_1,push_payload_0_0_0_0}}}}}}}}}}}}}}}}}}}};
  always @(posedge clk) begin
    if(popEvent_ready) begin
      tmp_ram_port0 <= ram[popPtr_value];
    end
  end

  always @(posedge clk) begin
    if(tmp_1) begin
      ram[pushPtr_value] <= tmp_ram_port;
    end
  end

  always @(*) begin
    tmp_1 = 1'b0;
    if(pushing) begin
      tmp_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 5'h1f);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + tmp_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 5'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 5'h1f);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + tmp_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 5'h0;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign pushing = (push_valid && push_ready);
  assign popping = (popEvent_valid && popEvent_ready);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign push_ready = (! full);
  assign popEvent_valid = ((! empty) && (! (tmp_popEvent_valid && (! full))));
  assign tmp_rData_0_0_0_0 = tmp_ram_port0;
  assign tmp_rData_0_0_0_0_1 = tmp_rData_0_0_0_0[1151 : 0];
  assign tmp_rData_0_0_0_0_2 = tmp_rData_0_0_0_0_1[383 : 0];
  assign tmp_rData_0_0_0_0_3 = tmp_rData_0_0_0_0_2[127 : 0];
  assign rData_0_0_0_0 = tmp_rData_0_0_0_0_3[7 : 0];
  assign rData_0_0_0_1 = tmp_rData_0_0_0_0_3[15 : 8];
  assign rData_0_0_0_2 = tmp_rData_0_0_0_0_3[23 : 16];
  assign rData_0_0_0_3 = tmp_rData_0_0_0_0_3[31 : 24];
  assign rData_0_0_0_4 = tmp_rData_0_0_0_0_3[39 : 32];
  assign rData_0_0_0_5 = tmp_rData_0_0_0_0_3[47 : 40];
  assign rData_0_0_0_6 = tmp_rData_0_0_0_0_3[55 : 48];
  assign rData_0_0_0_7 = tmp_rData_0_0_0_0_3[63 : 56];
  assign rData_0_0_0_8 = tmp_rData_0_0_0_0_3[71 : 64];
  assign rData_0_0_0_9 = tmp_rData_0_0_0_0_3[79 : 72];
  assign rData_0_0_0_10 = tmp_rData_0_0_0_0_3[87 : 80];
  assign rData_0_0_0_11 = tmp_rData_0_0_0_0_3[95 : 88];
  assign rData_0_0_0_12 = tmp_rData_0_0_0_0_3[103 : 96];
  assign rData_0_0_0_13 = tmp_rData_0_0_0_0_3[111 : 104];
  assign rData_0_0_0_14 = tmp_rData_0_0_0_0_3[119 : 112];
  assign rData_0_0_0_15 = tmp_rData_0_0_0_0_3[127 : 120];
  assign tmp_rData_0_0_1_0 = tmp_rData_0_0_0_0_2[255 : 128];
  assign rData_0_0_1_0 = tmp_rData_0_0_1_0[7 : 0];
  assign rData_0_0_1_1 = tmp_rData_0_0_1_0[15 : 8];
  assign rData_0_0_1_2 = tmp_rData_0_0_1_0[23 : 16];
  assign rData_0_0_1_3 = tmp_rData_0_0_1_0[31 : 24];
  assign rData_0_0_1_4 = tmp_rData_0_0_1_0[39 : 32];
  assign rData_0_0_1_5 = tmp_rData_0_0_1_0[47 : 40];
  assign rData_0_0_1_6 = tmp_rData_0_0_1_0[55 : 48];
  assign rData_0_0_1_7 = tmp_rData_0_0_1_0[63 : 56];
  assign rData_0_0_1_8 = tmp_rData_0_0_1_0[71 : 64];
  assign rData_0_0_1_9 = tmp_rData_0_0_1_0[79 : 72];
  assign rData_0_0_1_10 = tmp_rData_0_0_1_0[87 : 80];
  assign rData_0_0_1_11 = tmp_rData_0_0_1_0[95 : 88];
  assign rData_0_0_1_12 = tmp_rData_0_0_1_0[103 : 96];
  assign rData_0_0_1_13 = tmp_rData_0_0_1_0[111 : 104];
  assign rData_0_0_1_14 = tmp_rData_0_0_1_0[119 : 112];
  assign rData_0_0_1_15 = tmp_rData_0_0_1_0[127 : 120];
  assign tmp_rData_0_0_2_0 = tmp_rData_0_0_0_0_2[383 : 256];
  assign rData_0_0_2_0 = tmp_rData_0_0_2_0[7 : 0];
  assign rData_0_0_2_1 = tmp_rData_0_0_2_0[15 : 8];
  assign rData_0_0_2_2 = tmp_rData_0_0_2_0[23 : 16];
  assign rData_0_0_2_3 = tmp_rData_0_0_2_0[31 : 24];
  assign rData_0_0_2_4 = tmp_rData_0_0_2_0[39 : 32];
  assign rData_0_0_2_5 = tmp_rData_0_0_2_0[47 : 40];
  assign rData_0_0_2_6 = tmp_rData_0_0_2_0[55 : 48];
  assign rData_0_0_2_7 = tmp_rData_0_0_2_0[63 : 56];
  assign rData_0_0_2_8 = tmp_rData_0_0_2_0[71 : 64];
  assign rData_0_0_2_9 = tmp_rData_0_0_2_0[79 : 72];
  assign rData_0_0_2_10 = tmp_rData_0_0_2_0[87 : 80];
  assign rData_0_0_2_11 = tmp_rData_0_0_2_0[95 : 88];
  assign rData_0_0_2_12 = tmp_rData_0_0_2_0[103 : 96];
  assign rData_0_0_2_13 = tmp_rData_0_0_2_0[111 : 104];
  assign rData_0_0_2_14 = tmp_rData_0_0_2_0[119 : 112];
  assign rData_0_0_2_15 = tmp_rData_0_0_2_0[127 : 120];
  assign tmp_rData_0_1_0_0 = tmp_rData_0_0_0_0_1[767 : 384];
  assign tmp_rData_0_1_0_0_1 = tmp_rData_0_1_0_0[127 : 0];
  assign rData_0_1_0_0 = tmp_rData_0_1_0_0_1[7 : 0];
  assign rData_0_1_0_1 = tmp_rData_0_1_0_0_1[15 : 8];
  assign rData_0_1_0_2 = tmp_rData_0_1_0_0_1[23 : 16];
  assign rData_0_1_0_3 = tmp_rData_0_1_0_0_1[31 : 24];
  assign rData_0_1_0_4 = tmp_rData_0_1_0_0_1[39 : 32];
  assign rData_0_1_0_5 = tmp_rData_0_1_0_0_1[47 : 40];
  assign rData_0_1_0_6 = tmp_rData_0_1_0_0_1[55 : 48];
  assign rData_0_1_0_7 = tmp_rData_0_1_0_0_1[63 : 56];
  assign rData_0_1_0_8 = tmp_rData_0_1_0_0_1[71 : 64];
  assign rData_0_1_0_9 = tmp_rData_0_1_0_0_1[79 : 72];
  assign rData_0_1_0_10 = tmp_rData_0_1_0_0_1[87 : 80];
  assign rData_0_1_0_11 = tmp_rData_0_1_0_0_1[95 : 88];
  assign rData_0_1_0_12 = tmp_rData_0_1_0_0_1[103 : 96];
  assign rData_0_1_0_13 = tmp_rData_0_1_0_0_1[111 : 104];
  assign rData_0_1_0_14 = tmp_rData_0_1_0_0_1[119 : 112];
  assign rData_0_1_0_15 = tmp_rData_0_1_0_0_1[127 : 120];
  assign tmp_rData_0_1_1_0 = tmp_rData_0_1_0_0[255 : 128];
  assign rData_0_1_1_0 = tmp_rData_0_1_1_0[7 : 0];
  assign rData_0_1_1_1 = tmp_rData_0_1_1_0[15 : 8];
  assign rData_0_1_1_2 = tmp_rData_0_1_1_0[23 : 16];
  assign rData_0_1_1_3 = tmp_rData_0_1_1_0[31 : 24];
  assign rData_0_1_1_4 = tmp_rData_0_1_1_0[39 : 32];
  assign rData_0_1_1_5 = tmp_rData_0_1_1_0[47 : 40];
  assign rData_0_1_1_6 = tmp_rData_0_1_1_0[55 : 48];
  assign rData_0_1_1_7 = tmp_rData_0_1_1_0[63 : 56];
  assign rData_0_1_1_8 = tmp_rData_0_1_1_0[71 : 64];
  assign rData_0_1_1_9 = tmp_rData_0_1_1_0[79 : 72];
  assign rData_0_1_1_10 = tmp_rData_0_1_1_0[87 : 80];
  assign rData_0_1_1_11 = tmp_rData_0_1_1_0[95 : 88];
  assign rData_0_1_1_12 = tmp_rData_0_1_1_0[103 : 96];
  assign rData_0_1_1_13 = tmp_rData_0_1_1_0[111 : 104];
  assign rData_0_1_1_14 = tmp_rData_0_1_1_0[119 : 112];
  assign rData_0_1_1_15 = tmp_rData_0_1_1_0[127 : 120];
  assign tmp_rData_0_1_2_0 = tmp_rData_0_1_0_0[383 : 256];
  assign rData_0_1_2_0 = tmp_rData_0_1_2_0[7 : 0];
  assign rData_0_1_2_1 = tmp_rData_0_1_2_0[15 : 8];
  assign rData_0_1_2_2 = tmp_rData_0_1_2_0[23 : 16];
  assign rData_0_1_2_3 = tmp_rData_0_1_2_0[31 : 24];
  assign rData_0_1_2_4 = tmp_rData_0_1_2_0[39 : 32];
  assign rData_0_1_2_5 = tmp_rData_0_1_2_0[47 : 40];
  assign rData_0_1_2_6 = tmp_rData_0_1_2_0[55 : 48];
  assign rData_0_1_2_7 = tmp_rData_0_1_2_0[63 : 56];
  assign rData_0_1_2_8 = tmp_rData_0_1_2_0[71 : 64];
  assign rData_0_1_2_9 = tmp_rData_0_1_2_0[79 : 72];
  assign rData_0_1_2_10 = tmp_rData_0_1_2_0[87 : 80];
  assign rData_0_1_2_11 = tmp_rData_0_1_2_0[95 : 88];
  assign rData_0_1_2_12 = tmp_rData_0_1_2_0[103 : 96];
  assign rData_0_1_2_13 = tmp_rData_0_1_2_0[111 : 104];
  assign rData_0_1_2_14 = tmp_rData_0_1_2_0[119 : 112];
  assign rData_0_1_2_15 = tmp_rData_0_1_2_0[127 : 120];
  assign tmp_rData_0_2_0_0 = tmp_rData_0_0_0_0_1[1151 : 768];
  assign tmp_rData_0_2_0_0_1 = tmp_rData_0_2_0_0[127 : 0];
  assign rData_0_2_0_0 = tmp_rData_0_2_0_0_1[7 : 0];
  assign rData_0_2_0_1 = tmp_rData_0_2_0_0_1[15 : 8];
  assign rData_0_2_0_2 = tmp_rData_0_2_0_0_1[23 : 16];
  assign rData_0_2_0_3 = tmp_rData_0_2_0_0_1[31 : 24];
  assign rData_0_2_0_4 = tmp_rData_0_2_0_0_1[39 : 32];
  assign rData_0_2_0_5 = tmp_rData_0_2_0_0_1[47 : 40];
  assign rData_0_2_0_6 = tmp_rData_0_2_0_0_1[55 : 48];
  assign rData_0_2_0_7 = tmp_rData_0_2_0_0_1[63 : 56];
  assign rData_0_2_0_8 = tmp_rData_0_2_0_0_1[71 : 64];
  assign rData_0_2_0_9 = tmp_rData_0_2_0_0_1[79 : 72];
  assign rData_0_2_0_10 = tmp_rData_0_2_0_0_1[87 : 80];
  assign rData_0_2_0_11 = tmp_rData_0_2_0_0_1[95 : 88];
  assign rData_0_2_0_12 = tmp_rData_0_2_0_0_1[103 : 96];
  assign rData_0_2_0_13 = tmp_rData_0_2_0_0_1[111 : 104];
  assign rData_0_2_0_14 = tmp_rData_0_2_0_0_1[119 : 112];
  assign rData_0_2_0_15 = tmp_rData_0_2_0_0_1[127 : 120];
  assign tmp_rData_0_2_1_0 = tmp_rData_0_2_0_0[255 : 128];
  assign rData_0_2_1_0 = tmp_rData_0_2_1_0[7 : 0];
  assign rData_0_2_1_1 = tmp_rData_0_2_1_0[15 : 8];
  assign rData_0_2_1_2 = tmp_rData_0_2_1_0[23 : 16];
  assign rData_0_2_1_3 = tmp_rData_0_2_1_0[31 : 24];
  assign rData_0_2_1_4 = tmp_rData_0_2_1_0[39 : 32];
  assign rData_0_2_1_5 = tmp_rData_0_2_1_0[47 : 40];
  assign rData_0_2_1_6 = tmp_rData_0_2_1_0[55 : 48];
  assign rData_0_2_1_7 = tmp_rData_0_2_1_0[63 : 56];
  assign rData_0_2_1_8 = tmp_rData_0_2_1_0[71 : 64];
  assign rData_0_2_1_9 = tmp_rData_0_2_1_0[79 : 72];
  assign rData_0_2_1_10 = tmp_rData_0_2_1_0[87 : 80];
  assign rData_0_2_1_11 = tmp_rData_0_2_1_0[95 : 88];
  assign rData_0_2_1_12 = tmp_rData_0_2_1_0[103 : 96];
  assign rData_0_2_1_13 = tmp_rData_0_2_1_0[111 : 104];
  assign rData_0_2_1_14 = tmp_rData_0_2_1_0[119 : 112];
  assign rData_0_2_1_15 = tmp_rData_0_2_1_0[127 : 120];
  assign tmp_rData_0_2_2_0 = tmp_rData_0_2_0_0[383 : 256];
  assign rData_0_2_2_0 = tmp_rData_0_2_2_0[7 : 0];
  assign rData_0_2_2_1 = tmp_rData_0_2_2_0[15 : 8];
  assign rData_0_2_2_2 = tmp_rData_0_2_2_0[23 : 16];
  assign rData_0_2_2_3 = tmp_rData_0_2_2_0[31 : 24];
  assign rData_0_2_2_4 = tmp_rData_0_2_2_0[39 : 32];
  assign rData_0_2_2_5 = tmp_rData_0_2_2_0[47 : 40];
  assign rData_0_2_2_6 = tmp_rData_0_2_2_0[55 : 48];
  assign rData_0_2_2_7 = tmp_rData_0_2_2_0[63 : 56];
  assign rData_0_2_2_8 = tmp_rData_0_2_2_0[71 : 64];
  assign rData_0_2_2_9 = tmp_rData_0_2_2_0[79 : 72];
  assign rData_0_2_2_10 = tmp_rData_0_2_2_0[87 : 80];
  assign rData_0_2_2_11 = tmp_rData_0_2_2_0[95 : 88];
  assign rData_0_2_2_12 = tmp_rData_0_2_2_0[103 : 96];
  assign rData_0_2_2_13 = tmp_rData_0_2_2_0[111 : 104];
  assign rData_0_2_2_14 = tmp_rData_0_2_2_0[119 : 112];
  assign rData_0_2_2_15 = tmp_rData_0_2_2_0[127 : 120];
  assign tmp_rData_1_0_0_0 = tmp_rData_0_0_0_0[2303 : 1152];
  assign tmp_rData_1_0_0_0_1 = tmp_rData_1_0_0_0[383 : 0];
  assign tmp_rData_1_0_0_0_2 = tmp_rData_1_0_0_0_1[127 : 0];
  assign rData_1_0_0_0 = tmp_rData_1_0_0_0_2[7 : 0];
  assign rData_1_0_0_1 = tmp_rData_1_0_0_0_2[15 : 8];
  assign rData_1_0_0_2 = tmp_rData_1_0_0_0_2[23 : 16];
  assign rData_1_0_0_3 = tmp_rData_1_0_0_0_2[31 : 24];
  assign rData_1_0_0_4 = tmp_rData_1_0_0_0_2[39 : 32];
  assign rData_1_0_0_5 = tmp_rData_1_0_0_0_2[47 : 40];
  assign rData_1_0_0_6 = tmp_rData_1_0_0_0_2[55 : 48];
  assign rData_1_0_0_7 = tmp_rData_1_0_0_0_2[63 : 56];
  assign rData_1_0_0_8 = tmp_rData_1_0_0_0_2[71 : 64];
  assign rData_1_0_0_9 = tmp_rData_1_0_0_0_2[79 : 72];
  assign rData_1_0_0_10 = tmp_rData_1_0_0_0_2[87 : 80];
  assign rData_1_0_0_11 = tmp_rData_1_0_0_0_2[95 : 88];
  assign rData_1_0_0_12 = tmp_rData_1_0_0_0_2[103 : 96];
  assign rData_1_0_0_13 = tmp_rData_1_0_0_0_2[111 : 104];
  assign rData_1_0_0_14 = tmp_rData_1_0_0_0_2[119 : 112];
  assign rData_1_0_0_15 = tmp_rData_1_0_0_0_2[127 : 120];
  assign tmp_rData_1_0_1_0 = tmp_rData_1_0_0_0_1[255 : 128];
  assign rData_1_0_1_0 = tmp_rData_1_0_1_0[7 : 0];
  assign rData_1_0_1_1 = tmp_rData_1_0_1_0[15 : 8];
  assign rData_1_0_1_2 = tmp_rData_1_0_1_0[23 : 16];
  assign rData_1_0_1_3 = tmp_rData_1_0_1_0[31 : 24];
  assign rData_1_0_1_4 = tmp_rData_1_0_1_0[39 : 32];
  assign rData_1_0_1_5 = tmp_rData_1_0_1_0[47 : 40];
  assign rData_1_0_1_6 = tmp_rData_1_0_1_0[55 : 48];
  assign rData_1_0_1_7 = tmp_rData_1_0_1_0[63 : 56];
  assign rData_1_0_1_8 = tmp_rData_1_0_1_0[71 : 64];
  assign rData_1_0_1_9 = tmp_rData_1_0_1_0[79 : 72];
  assign rData_1_0_1_10 = tmp_rData_1_0_1_0[87 : 80];
  assign rData_1_0_1_11 = tmp_rData_1_0_1_0[95 : 88];
  assign rData_1_0_1_12 = tmp_rData_1_0_1_0[103 : 96];
  assign rData_1_0_1_13 = tmp_rData_1_0_1_0[111 : 104];
  assign rData_1_0_1_14 = tmp_rData_1_0_1_0[119 : 112];
  assign rData_1_0_1_15 = tmp_rData_1_0_1_0[127 : 120];
  assign tmp_rData_1_0_2_0 = tmp_rData_1_0_0_0_1[383 : 256];
  assign rData_1_0_2_0 = tmp_rData_1_0_2_0[7 : 0];
  assign rData_1_0_2_1 = tmp_rData_1_0_2_0[15 : 8];
  assign rData_1_0_2_2 = tmp_rData_1_0_2_0[23 : 16];
  assign rData_1_0_2_3 = tmp_rData_1_0_2_0[31 : 24];
  assign rData_1_0_2_4 = tmp_rData_1_0_2_0[39 : 32];
  assign rData_1_0_2_5 = tmp_rData_1_0_2_0[47 : 40];
  assign rData_1_0_2_6 = tmp_rData_1_0_2_0[55 : 48];
  assign rData_1_0_2_7 = tmp_rData_1_0_2_0[63 : 56];
  assign rData_1_0_2_8 = tmp_rData_1_0_2_0[71 : 64];
  assign rData_1_0_2_9 = tmp_rData_1_0_2_0[79 : 72];
  assign rData_1_0_2_10 = tmp_rData_1_0_2_0[87 : 80];
  assign rData_1_0_2_11 = tmp_rData_1_0_2_0[95 : 88];
  assign rData_1_0_2_12 = tmp_rData_1_0_2_0[103 : 96];
  assign rData_1_0_2_13 = tmp_rData_1_0_2_0[111 : 104];
  assign rData_1_0_2_14 = tmp_rData_1_0_2_0[119 : 112];
  assign rData_1_0_2_15 = tmp_rData_1_0_2_0[127 : 120];
  assign tmp_rData_1_1_0_0 = tmp_rData_1_0_0_0[767 : 384];
  assign tmp_rData_1_1_0_0_1 = tmp_rData_1_1_0_0[127 : 0];
  assign rData_1_1_0_0 = tmp_rData_1_1_0_0_1[7 : 0];
  assign rData_1_1_0_1 = tmp_rData_1_1_0_0_1[15 : 8];
  assign rData_1_1_0_2 = tmp_rData_1_1_0_0_1[23 : 16];
  assign rData_1_1_0_3 = tmp_rData_1_1_0_0_1[31 : 24];
  assign rData_1_1_0_4 = tmp_rData_1_1_0_0_1[39 : 32];
  assign rData_1_1_0_5 = tmp_rData_1_1_0_0_1[47 : 40];
  assign rData_1_1_0_6 = tmp_rData_1_1_0_0_1[55 : 48];
  assign rData_1_1_0_7 = tmp_rData_1_1_0_0_1[63 : 56];
  assign rData_1_1_0_8 = tmp_rData_1_1_0_0_1[71 : 64];
  assign rData_1_1_0_9 = tmp_rData_1_1_0_0_1[79 : 72];
  assign rData_1_1_0_10 = tmp_rData_1_1_0_0_1[87 : 80];
  assign rData_1_1_0_11 = tmp_rData_1_1_0_0_1[95 : 88];
  assign rData_1_1_0_12 = tmp_rData_1_1_0_0_1[103 : 96];
  assign rData_1_1_0_13 = tmp_rData_1_1_0_0_1[111 : 104];
  assign rData_1_1_0_14 = tmp_rData_1_1_0_0_1[119 : 112];
  assign rData_1_1_0_15 = tmp_rData_1_1_0_0_1[127 : 120];
  assign tmp_rData_1_1_1_0 = tmp_rData_1_1_0_0[255 : 128];
  assign rData_1_1_1_0 = tmp_rData_1_1_1_0[7 : 0];
  assign rData_1_1_1_1 = tmp_rData_1_1_1_0[15 : 8];
  assign rData_1_1_1_2 = tmp_rData_1_1_1_0[23 : 16];
  assign rData_1_1_1_3 = tmp_rData_1_1_1_0[31 : 24];
  assign rData_1_1_1_4 = tmp_rData_1_1_1_0[39 : 32];
  assign rData_1_1_1_5 = tmp_rData_1_1_1_0[47 : 40];
  assign rData_1_1_1_6 = tmp_rData_1_1_1_0[55 : 48];
  assign rData_1_1_1_7 = tmp_rData_1_1_1_0[63 : 56];
  assign rData_1_1_1_8 = tmp_rData_1_1_1_0[71 : 64];
  assign rData_1_1_1_9 = tmp_rData_1_1_1_0[79 : 72];
  assign rData_1_1_1_10 = tmp_rData_1_1_1_0[87 : 80];
  assign rData_1_1_1_11 = tmp_rData_1_1_1_0[95 : 88];
  assign rData_1_1_1_12 = tmp_rData_1_1_1_0[103 : 96];
  assign rData_1_1_1_13 = tmp_rData_1_1_1_0[111 : 104];
  assign rData_1_1_1_14 = tmp_rData_1_1_1_0[119 : 112];
  assign rData_1_1_1_15 = tmp_rData_1_1_1_0[127 : 120];
  assign tmp_rData_1_1_2_0 = tmp_rData_1_1_0_0[383 : 256];
  assign rData_1_1_2_0 = tmp_rData_1_1_2_0[7 : 0];
  assign rData_1_1_2_1 = tmp_rData_1_1_2_0[15 : 8];
  assign rData_1_1_2_2 = tmp_rData_1_1_2_0[23 : 16];
  assign rData_1_1_2_3 = tmp_rData_1_1_2_0[31 : 24];
  assign rData_1_1_2_4 = tmp_rData_1_1_2_0[39 : 32];
  assign rData_1_1_2_5 = tmp_rData_1_1_2_0[47 : 40];
  assign rData_1_1_2_6 = tmp_rData_1_1_2_0[55 : 48];
  assign rData_1_1_2_7 = tmp_rData_1_1_2_0[63 : 56];
  assign rData_1_1_2_8 = tmp_rData_1_1_2_0[71 : 64];
  assign rData_1_1_2_9 = tmp_rData_1_1_2_0[79 : 72];
  assign rData_1_1_2_10 = tmp_rData_1_1_2_0[87 : 80];
  assign rData_1_1_2_11 = tmp_rData_1_1_2_0[95 : 88];
  assign rData_1_1_2_12 = tmp_rData_1_1_2_0[103 : 96];
  assign rData_1_1_2_13 = tmp_rData_1_1_2_0[111 : 104];
  assign rData_1_1_2_14 = tmp_rData_1_1_2_0[119 : 112];
  assign rData_1_1_2_15 = tmp_rData_1_1_2_0[127 : 120];
  assign tmp_rData_1_2_0_0 = tmp_rData_1_0_0_0[1151 : 768];
  assign tmp_rData_1_2_0_0_1 = tmp_rData_1_2_0_0[127 : 0];
  assign rData_1_2_0_0 = tmp_rData_1_2_0_0_1[7 : 0];
  assign rData_1_2_0_1 = tmp_rData_1_2_0_0_1[15 : 8];
  assign rData_1_2_0_2 = tmp_rData_1_2_0_0_1[23 : 16];
  assign rData_1_2_0_3 = tmp_rData_1_2_0_0_1[31 : 24];
  assign rData_1_2_0_4 = tmp_rData_1_2_0_0_1[39 : 32];
  assign rData_1_2_0_5 = tmp_rData_1_2_0_0_1[47 : 40];
  assign rData_1_2_0_6 = tmp_rData_1_2_0_0_1[55 : 48];
  assign rData_1_2_0_7 = tmp_rData_1_2_0_0_1[63 : 56];
  assign rData_1_2_0_8 = tmp_rData_1_2_0_0_1[71 : 64];
  assign rData_1_2_0_9 = tmp_rData_1_2_0_0_1[79 : 72];
  assign rData_1_2_0_10 = tmp_rData_1_2_0_0_1[87 : 80];
  assign rData_1_2_0_11 = tmp_rData_1_2_0_0_1[95 : 88];
  assign rData_1_2_0_12 = tmp_rData_1_2_0_0_1[103 : 96];
  assign rData_1_2_0_13 = tmp_rData_1_2_0_0_1[111 : 104];
  assign rData_1_2_0_14 = tmp_rData_1_2_0_0_1[119 : 112];
  assign rData_1_2_0_15 = tmp_rData_1_2_0_0_1[127 : 120];
  assign tmp_rData_1_2_1_0 = tmp_rData_1_2_0_0[255 : 128];
  assign rData_1_2_1_0 = tmp_rData_1_2_1_0[7 : 0];
  assign rData_1_2_1_1 = tmp_rData_1_2_1_0[15 : 8];
  assign rData_1_2_1_2 = tmp_rData_1_2_1_0[23 : 16];
  assign rData_1_2_1_3 = tmp_rData_1_2_1_0[31 : 24];
  assign rData_1_2_1_4 = tmp_rData_1_2_1_0[39 : 32];
  assign rData_1_2_1_5 = tmp_rData_1_2_1_0[47 : 40];
  assign rData_1_2_1_6 = tmp_rData_1_2_1_0[55 : 48];
  assign rData_1_2_1_7 = tmp_rData_1_2_1_0[63 : 56];
  assign rData_1_2_1_8 = tmp_rData_1_2_1_0[71 : 64];
  assign rData_1_2_1_9 = tmp_rData_1_2_1_0[79 : 72];
  assign rData_1_2_1_10 = tmp_rData_1_2_1_0[87 : 80];
  assign rData_1_2_1_11 = tmp_rData_1_2_1_0[95 : 88];
  assign rData_1_2_1_12 = tmp_rData_1_2_1_0[103 : 96];
  assign rData_1_2_1_13 = tmp_rData_1_2_1_0[111 : 104];
  assign rData_1_2_1_14 = tmp_rData_1_2_1_0[119 : 112];
  assign rData_1_2_1_15 = tmp_rData_1_2_1_0[127 : 120];
  assign tmp_rData_1_2_2_0 = tmp_rData_1_2_0_0[383 : 256];
  assign rData_1_2_2_0 = tmp_rData_1_2_2_0[7 : 0];
  assign rData_1_2_2_1 = tmp_rData_1_2_2_0[15 : 8];
  assign rData_1_2_2_2 = tmp_rData_1_2_2_0[23 : 16];
  assign rData_1_2_2_3 = tmp_rData_1_2_2_0[31 : 24];
  assign rData_1_2_2_4 = tmp_rData_1_2_2_0[39 : 32];
  assign rData_1_2_2_5 = tmp_rData_1_2_2_0[47 : 40];
  assign rData_1_2_2_6 = tmp_rData_1_2_2_0[55 : 48];
  assign rData_1_2_2_7 = tmp_rData_1_2_2_0[63 : 56];
  assign rData_1_2_2_8 = tmp_rData_1_2_2_0[71 : 64];
  assign rData_1_2_2_9 = tmp_rData_1_2_2_0[79 : 72];
  assign rData_1_2_2_10 = tmp_rData_1_2_2_0[87 : 80];
  assign rData_1_2_2_11 = tmp_rData_1_2_2_0[95 : 88];
  assign rData_1_2_2_12 = tmp_rData_1_2_2_0[103 : 96];
  assign rData_1_2_2_13 = tmp_rData_1_2_2_0[111 : 104];
  assign rData_1_2_2_14 = tmp_rData_1_2_2_0[119 : 112];
  assign rData_1_2_2_15 = tmp_rData_1_2_2_0[127 : 120];
  always @(*) begin
    popEvent_ready = pop_ready;
    if(when_StreamFifoHighPerf_l38) begin
      popEvent_ready = 1'b1;
    end
  end

  assign when_StreamFifoHighPerf_l38 = (! rValid);
  assign pop_valid = rValid;
  assign pop_payload_0_0_0_0 = rData_0_0_0_0;
  assign pop_payload_0_0_0_1 = rData_0_0_0_1;
  assign pop_payload_0_0_0_2 = rData_0_0_0_2;
  assign pop_payload_0_0_0_3 = rData_0_0_0_3;
  assign pop_payload_0_0_0_4 = rData_0_0_0_4;
  assign pop_payload_0_0_0_5 = rData_0_0_0_5;
  assign pop_payload_0_0_0_6 = rData_0_0_0_6;
  assign pop_payload_0_0_0_7 = rData_0_0_0_7;
  assign pop_payload_0_0_0_8 = rData_0_0_0_8;
  assign pop_payload_0_0_0_9 = rData_0_0_0_9;
  assign pop_payload_0_0_0_10 = rData_0_0_0_10;
  assign pop_payload_0_0_0_11 = rData_0_0_0_11;
  assign pop_payload_0_0_0_12 = rData_0_0_0_12;
  assign pop_payload_0_0_0_13 = rData_0_0_0_13;
  assign pop_payload_0_0_0_14 = rData_0_0_0_14;
  assign pop_payload_0_0_0_15 = rData_0_0_0_15;
  assign pop_payload_0_0_1_0 = rData_0_0_1_0;
  assign pop_payload_0_0_1_1 = rData_0_0_1_1;
  assign pop_payload_0_0_1_2 = rData_0_0_1_2;
  assign pop_payload_0_0_1_3 = rData_0_0_1_3;
  assign pop_payload_0_0_1_4 = rData_0_0_1_4;
  assign pop_payload_0_0_1_5 = rData_0_0_1_5;
  assign pop_payload_0_0_1_6 = rData_0_0_1_6;
  assign pop_payload_0_0_1_7 = rData_0_0_1_7;
  assign pop_payload_0_0_1_8 = rData_0_0_1_8;
  assign pop_payload_0_0_1_9 = rData_0_0_1_9;
  assign pop_payload_0_0_1_10 = rData_0_0_1_10;
  assign pop_payload_0_0_1_11 = rData_0_0_1_11;
  assign pop_payload_0_0_1_12 = rData_0_0_1_12;
  assign pop_payload_0_0_1_13 = rData_0_0_1_13;
  assign pop_payload_0_0_1_14 = rData_0_0_1_14;
  assign pop_payload_0_0_1_15 = rData_0_0_1_15;
  assign pop_payload_0_0_2_0 = rData_0_0_2_0;
  assign pop_payload_0_0_2_1 = rData_0_0_2_1;
  assign pop_payload_0_0_2_2 = rData_0_0_2_2;
  assign pop_payload_0_0_2_3 = rData_0_0_2_3;
  assign pop_payload_0_0_2_4 = rData_0_0_2_4;
  assign pop_payload_0_0_2_5 = rData_0_0_2_5;
  assign pop_payload_0_0_2_6 = rData_0_0_2_6;
  assign pop_payload_0_0_2_7 = rData_0_0_2_7;
  assign pop_payload_0_0_2_8 = rData_0_0_2_8;
  assign pop_payload_0_0_2_9 = rData_0_0_2_9;
  assign pop_payload_0_0_2_10 = rData_0_0_2_10;
  assign pop_payload_0_0_2_11 = rData_0_0_2_11;
  assign pop_payload_0_0_2_12 = rData_0_0_2_12;
  assign pop_payload_0_0_2_13 = rData_0_0_2_13;
  assign pop_payload_0_0_2_14 = rData_0_0_2_14;
  assign pop_payload_0_0_2_15 = rData_0_0_2_15;
  assign pop_payload_0_1_0_0 = rData_0_1_0_0;
  assign pop_payload_0_1_0_1 = rData_0_1_0_1;
  assign pop_payload_0_1_0_2 = rData_0_1_0_2;
  assign pop_payload_0_1_0_3 = rData_0_1_0_3;
  assign pop_payload_0_1_0_4 = rData_0_1_0_4;
  assign pop_payload_0_1_0_5 = rData_0_1_0_5;
  assign pop_payload_0_1_0_6 = rData_0_1_0_6;
  assign pop_payload_0_1_0_7 = rData_0_1_0_7;
  assign pop_payload_0_1_0_8 = rData_0_1_0_8;
  assign pop_payload_0_1_0_9 = rData_0_1_0_9;
  assign pop_payload_0_1_0_10 = rData_0_1_0_10;
  assign pop_payload_0_1_0_11 = rData_0_1_0_11;
  assign pop_payload_0_1_0_12 = rData_0_1_0_12;
  assign pop_payload_0_1_0_13 = rData_0_1_0_13;
  assign pop_payload_0_1_0_14 = rData_0_1_0_14;
  assign pop_payload_0_1_0_15 = rData_0_1_0_15;
  assign pop_payload_0_1_1_0 = rData_0_1_1_0;
  assign pop_payload_0_1_1_1 = rData_0_1_1_1;
  assign pop_payload_0_1_1_2 = rData_0_1_1_2;
  assign pop_payload_0_1_1_3 = rData_0_1_1_3;
  assign pop_payload_0_1_1_4 = rData_0_1_1_4;
  assign pop_payload_0_1_1_5 = rData_0_1_1_5;
  assign pop_payload_0_1_1_6 = rData_0_1_1_6;
  assign pop_payload_0_1_1_7 = rData_0_1_1_7;
  assign pop_payload_0_1_1_8 = rData_0_1_1_8;
  assign pop_payload_0_1_1_9 = rData_0_1_1_9;
  assign pop_payload_0_1_1_10 = rData_0_1_1_10;
  assign pop_payload_0_1_1_11 = rData_0_1_1_11;
  assign pop_payload_0_1_1_12 = rData_0_1_1_12;
  assign pop_payload_0_1_1_13 = rData_0_1_1_13;
  assign pop_payload_0_1_1_14 = rData_0_1_1_14;
  assign pop_payload_0_1_1_15 = rData_0_1_1_15;
  assign pop_payload_0_1_2_0 = rData_0_1_2_0;
  assign pop_payload_0_1_2_1 = rData_0_1_2_1;
  assign pop_payload_0_1_2_2 = rData_0_1_2_2;
  assign pop_payload_0_1_2_3 = rData_0_1_2_3;
  assign pop_payload_0_1_2_4 = rData_0_1_2_4;
  assign pop_payload_0_1_2_5 = rData_0_1_2_5;
  assign pop_payload_0_1_2_6 = rData_0_1_2_6;
  assign pop_payload_0_1_2_7 = rData_0_1_2_7;
  assign pop_payload_0_1_2_8 = rData_0_1_2_8;
  assign pop_payload_0_1_2_9 = rData_0_1_2_9;
  assign pop_payload_0_1_2_10 = rData_0_1_2_10;
  assign pop_payload_0_1_2_11 = rData_0_1_2_11;
  assign pop_payload_0_1_2_12 = rData_0_1_2_12;
  assign pop_payload_0_1_2_13 = rData_0_1_2_13;
  assign pop_payload_0_1_2_14 = rData_0_1_2_14;
  assign pop_payload_0_1_2_15 = rData_0_1_2_15;
  assign pop_payload_0_2_0_0 = rData_0_2_0_0;
  assign pop_payload_0_2_0_1 = rData_0_2_0_1;
  assign pop_payload_0_2_0_2 = rData_0_2_0_2;
  assign pop_payload_0_2_0_3 = rData_0_2_0_3;
  assign pop_payload_0_2_0_4 = rData_0_2_0_4;
  assign pop_payload_0_2_0_5 = rData_0_2_0_5;
  assign pop_payload_0_2_0_6 = rData_0_2_0_6;
  assign pop_payload_0_2_0_7 = rData_0_2_0_7;
  assign pop_payload_0_2_0_8 = rData_0_2_0_8;
  assign pop_payload_0_2_0_9 = rData_0_2_0_9;
  assign pop_payload_0_2_0_10 = rData_0_2_0_10;
  assign pop_payload_0_2_0_11 = rData_0_2_0_11;
  assign pop_payload_0_2_0_12 = rData_0_2_0_12;
  assign pop_payload_0_2_0_13 = rData_0_2_0_13;
  assign pop_payload_0_2_0_14 = rData_0_2_0_14;
  assign pop_payload_0_2_0_15 = rData_0_2_0_15;
  assign pop_payload_0_2_1_0 = rData_0_2_1_0;
  assign pop_payload_0_2_1_1 = rData_0_2_1_1;
  assign pop_payload_0_2_1_2 = rData_0_2_1_2;
  assign pop_payload_0_2_1_3 = rData_0_2_1_3;
  assign pop_payload_0_2_1_4 = rData_0_2_1_4;
  assign pop_payload_0_2_1_5 = rData_0_2_1_5;
  assign pop_payload_0_2_1_6 = rData_0_2_1_6;
  assign pop_payload_0_2_1_7 = rData_0_2_1_7;
  assign pop_payload_0_2_1_8 = rData_0_2_1_8;
  assign pop_payload_0_2_1_9 = rData_0_2_1_9;
  assign pop_payload_0_2_1_10 = rData_0_2_1_10;
  assign pop_payload_0_2_1_11 = rData_0_2_1_11;
  assign pop_payload_0_2_1_12 = rData_0_2_1_12;
  assign pop_payload_0_2_1_13 = rData_0_2_1_13;
  assign pop_payload_0_2_1_14 = rData_0_2_1_14;
  assign pop_payload_0_2_1_15 = rData_0_2_1_15;
  assign pop_payload_0_2_2_0 = rData_0_2_2_0;
  assign pop_payload_0_2_2_1 = rData_0_2_2_1;
  assign pop_payload_0_2_2_2 = rData_0_2_2_2;
  assign pop_payload_0_2_2_3 = rData_0_2_2_3;
  assign pop_payload_0_2_2_4 = rData_0_2_2_4;
  assign pop_payload_0_2_2_5 = rData_0_2_2_5;
  assign pop_payload_0_2_2_6 = rData_0_2_2_6;
  assign pop_payload_0_2_2_7 = rData_0_2_2_7;
  assign pop_payload_0_2_2_8 = rData_0_2_2_8;
  assign pop_payload_0_2_2_9 = rData_0_2_2_9;
  assign pop_payload_0_2_2_10 = rData_0_2_2_10;
  assign pop_payload_0_2_2_11 = rData_0_2_2_11;
  assign pop_payload_0_2_2_12 = rData_0_2_2_12;
  assign pop_payload_0_2_2_13 = rData_0_2_2_13;
  assign pop_payload_0_2_2_14 = rData_0_2_2_14;
  assign pop_payload_0_2_2_15 = rData_0_2_2_15;
  assign pop_payload_1_0_0_0 = rData_1_0_0_0;
  assign pop_payload_1_0_0_1 = rData_1_0_0_1;
  assign pop_payload_1_0_0_2 = rData_1_0_0_2;
  assign pop_payload_1_0_0_3 = rData_1_0_0_3;
  assign pop_payload_1_0_0_4 = rData_1_0_0_4;
  assign pop_payload_1_0_0_5 = rData_1_0_0_5;
  assign pop_payload_1_0_0_6 = rData_1_0_0_6;
  assign pop_payload_1_0_0_7 = rData_1_0_0_7;
  assign pop_payload_1_0_0_8 = rData_1_0_0_8;
  assign pop_payload_1_0_0_9 = rData_1_0_0_9;
  assign pop_payload_1_0_0_10 = rData_1_0_0_10;
  assign pop_payload_1_0_0_11 = rData_1_0_0_11;
  assign pop_payload_1_0_0_12 = rData_1_0_0_12;
  assign pop_payload_1_0_0_13 = rData_1_0_0_13;
  assign pop_payload_1_0_0_14 = rData_1_0_0_14;
  assign pop_payload_1_0_0_15 = rData_1_0_0_15;
  assign pop_payload_1_0_1_0 = rData_1_0_1_0;
  assign pop_payload_1_0_1_1 = rData_1_0_1_1;
  assign pop_payload_1_0_1_2 = rData_1_0_1_2;
  assign pop_payload_1_0_1_3 = rData_1_0_1_3;
  assign pop_payload_1_0_1_4 = rData_1_0_1_4;
  assign pop_payload_1_0_1_5 = rData_1_0_1_5;
  assign pop_payload_1_0_1_6 = rData_1_0_1_6;
  assign pop_payload_1_0_1_7 = rData_1_0_1_7;
  assign pop_payload_1_0_1_8 = rData_1_0_1_8;
  assign pop_payload_1_0_1_9 = rData_1_0_1_9;
  assign pop_payload_1_0_1_10 = rData_1_0_1_10;
  assign pop_payload_1_0_1_11 = rData_1_0_1_11;
  assign pop_payload_1_0_1_12 = rData_1_0_1_12;
  assign pop_payload_1_0_1_13 = rData_1_0_1_13;
  assign pop_payload_1_0_1_14 = rData_1_0_1_14;
  assign pop_payload_1_0_1_15 = rData_1_0_1_15;
  assign pop_payload_1_0_2_0 = rData_1_0_2_0;
  assign pop_payload_1_0_2_1 = rData_1_0_2_1;
  assign pop_payload_1_0_2_2 = rData_1_0_2_2;
  assign pop_payload_1_0_2_3 = rData_1_0_2_3;
  assign pop_payload_1_0_2_4 = rData_1_0_2_4;
  assign pop_payload_1_0_2_5 = rData_1_0_2_5;
  assign pop_payload_1_0_2_6 = rData_1_0_2_6;
  assign pop_payload_1_0_2_7 = rData_1_0_2_7;
  assign pop_payload_1_0_2_8 = rData_1_0_2_8;
  assign pop_payload_1_0_2_9 = rData_1_0_2_9;
  assign pop_payload_1_0_2_10 = rData_1_0_2_10;
  assign pop_payload_1_0_2_11 = rData_1_0_2_11;
  assign pop_payload_1_0_2_12 = rData_1_0_2_12;
  assign pop_payload_1_0_2_13 = rData_1_0_2_13;
  assign pop_payload_1_0_2_14 = rData_1_0_2_14;
  assign pop_payload_1_0_2_15 = rData_1_0_2_15;
  assign pop_payload_1_1_0_0 = rData_1_1_0_0;
  assign pop_payload_1_1_0_1 = rData_1_1_0_1;
  assign pop_payload_1_1_0_2 = rData_1_1_0_2;
  assign pop_payload_1_1_0_3 = rData_1_1_0_3;
  assign pop_payload_1_1_0_4 = rData_1_1_0_4;
  assign pop_payload_1_1_0_5 = rData_1_1_0_5;
  assign pop_payload_1_1_0_6 = rData_1_1_0_6;
  assign pop_payload_1_1_0_7 = rData_1_1_0_7;
  assign pop_payload_1_1_0_8 = rData_1_1_0_8;
  assign pop_payload_1_1_0_9 = rData_1_1_0_9;
  assign pop_payload_1_1_0_10 = rData_1_1_0_10;
  assign pop_payload_1_1_0_11 = rData_1_1_0_11;
  assign pop_payload_1_1_0_12 = rData_1_1_0_12;
  assign pop_payload_1_1_0_13 = rData_1_1_0_13;
  assign pop_payload_1_1_0_14 = rData_1_1_0_14;
  assign pop_payload_1_1_0_15 = rData_1_1_0_15;
  assign pop_payload_1_1_1_0 = rData_1_1_1_0;
  assign pop_payload_1_1_1_1 = rData_1_1_1_1;
  assign pop_payload_1_1_1_2 = rData_1_1_1_2;
  assign pop_payload_1_1_1_3 = rData_1_1_1_3;
  assign pop_payload_1_1_1_4 = rData_1_1_1_4;
  assign pop_payload_1_1_1_5 = rData_1_1_1_5;
  assign pop_payload_1_1_1_6 = rData_1_1_1_6;
  assign pop_payload_1_1_1_7 = rData_1_1_1_7;
  assign pop_payload_1_1_1_8 = rData_1_1_1_8;
  assign pop_payload_1_1_1_9 = rData_1_1_1_9;
  assign pop_payload_1_1_1_10 = rData_1_1_1_10;
  assign pop_payload_1_1_1_11 = rData_1_1_1_11;
  assign pop_payload_1_1_1_12 = rData_1_1_1_12;
  assign pop_payload_1_1_1_13 = rData_1_1_1_13;
  assign pop_payload_1_1_1_14 = rData_1_1_1_14;
  assign pop_payload_1_1_1_15 = rData_1_1_1_15;
  assign pop_payload_1_1_2_0 = rData_1_1_2_0;
  assign pop_payload_1_1_2_1 = rData_1_1_2_1;
  assign pop_payload_1_1_2_2 = rData_1_1_2_2;
  assign pop_payload_1_1_2_3 = rData_1_1_2_3;
  assign pop_payload_1_1_2_4 = rData_1_1_2_4;
  assign pop_payload_1_1_2_5 = rData_1_1_2_5;
  assign pop_payload_1_1_2_6 = rData_1_1_2_6;
  assign pop_payload_1_1_2_7 = rData_1_1_2_7;
  assign pop_payload_1_1_2_8 = rData_1_1_2_8;
  assign pop_payload_1_1_2_9 = rData_1_1_2_9;
  assign pop_payload_1_1_2_10 = rData_1_1_2_10;
  assign pop_payload_1_1_2_11 = rData_1_1_2_11;
  assign pop_payload_1_1_2_12 = rData_1_1_2_12;
  assign pop_payload_1_1_2_13 = rData_1_1_2_13;
  assign pop_payload_1_1_2_14 = rData_1_1_2_14;
  assign pop_payload_1_1_2_15 = rData_1_1_2_15;
  assign pop_payload_1_2_0_0 = rData_1_2_0_0;
  assign pop_payload_1_2_0_1 = rData_1_2_0_1;
  assign pop_payload_1_2_0_2 = rData_1_2_0_2;
  assign pop_payload_1_2_0_3 = rData_1_2_0_3;
  assign pop_payload_1_2_0_4 = rData_1_2_0_4;
  assign pop_payload_1_2_0_5 = rData_1_2_0_5;
  assign pop_payload_1_2_0_6 = rData_1_2_0_6;
  assign pop_payload_1_2_0_7 = rData_1_2_0_7;
  assign pop_payload_1_2_0_8 = rData_1_2_0_8;
  assign pop_payload_1_2_0_9 = rData_1_2_0_9;
  assign pop_payload_1_2_0_10 = rData_1_2_0_10;
  assign pop_payload_1_2_0_11 = rData_1_2_0_11;
  assign pop_payload_1_2_0_12 = rData_1_2_0_12;
  assign pop_payload_1_2_0_13 = rData_1_2_0_13;
  assign pop_payload_1_2_0_14 = rData_1_2_0_14;
  assign pop_payload_1_2_0_15 = rData_1_2_0_15;
  assign pop_payload_1_2_1_0 = rData_1_2_1_0;
  assign pop_payload_1_2_1_1 = rData_1_2_1_1;
  assign pop_payload_1_2_1_2 = rData_1_2_1_2;
  assign pop_payload_1_2_1_3 = rData_1_2_1_3;
  assign pop_payload_1_2_1_4 = rData_1_2_1_4;
  assign pop_payload_1_2_1_5 = rData_1_2_1_5;
  assign pop_payload_1_2_1_6 = rData_1_2_1_6;
  assign pop_payload_1_2_1_7 = rData_1_2_1_7;
  assign pop_payload_1_2_1_8 = rData_1_2_1_8;
  assign pop_payload_1_2_1_9 = rData_1_2_1_9;
  assign pop_payload_1_2_1_10 = rData_1_2_1_10;
  assign pop_payload_1_2_1_11 = rData_1_2_1_11;
  assign pop_payload_1_2_1_12 = rData_1_2_1_12;
  assign pop_payload_1_2_1_13 = rData_1_2_1_13;
  assign pop_payload_1_2_1_14 = rData_1_2_1_14;
  assign pop_payload_1_2_1_15 = rData_1_2_1_15;
  assign pop_payload_1_2_2_0 = rData_1_2_2_0;
  assign pop_payload_1_2_2_1 = rData_1_2_2_1;
  assign pop_payload_1_2_2_2 = rData_1_2_2_2;
  assign pop_payload_1_2_2_3 = rData_1_2_2_3;
  assign pop_payload_1_2_2_4 = rData_1_2_2_4;
  assign pop_payload_1_2_2_5 = rData_1_2_2_5;
  assign pop_payload_1_2_2_6 = rData_1_2_2_6;
  assign pop_payload_1_2_2_7 = rData_1_2_2_7;
  assign pop_payload_1_2_2_8 = rData_1_2_2_8;
  assign pop_payload_1_2_2_9 = rData_1_2_2_9;
  assign pop_payload_1_2_2_10 = rData_1_2_2_10;
  assign pop_payload_1_2_2_11 = rData_1_2_2_11;
  assign pop_payload_1_2_2_12 = rData_1_2_2_12;
  assign pop_payload_1_2_2_13 = rData_1_2_2_13;
  assign pop_payload_1_2_2_14 = rData_1_2_2_14;
  assign pop_payload_1_2_2_15 = rData_1_2_2_15;
  assign when_StreamFifoHighPerf_l42 = (pushing != popping);
  always @(posedge clk) begin
    if(reset) begin
      pushPtr_value <= 5'h0;
      popPtr_value <= 5'h0;
      risingOccupancy <= 1'b0;
      tmp_popEvent_valid <= 1'b0;
      rValid <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      tmp_popEvent_valid <= (popPtr_valueNext == pushPtr_value);
      if(popEvent_ready) begin
        rValid <= popEvent_valid;
      end
      if(when_StreamFifoHighPerf_l42) begin
        risingOccupancy <= pushing;
      end
      if(flush) begin
        rValid <= 1'b0;
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

//SInt48fixTo7_0_ROUNDTOINF replaced by SInt48fixTo7_0_ROUNDTOINF

//AMultB replaced by AMultB

module SInt48fixTo7_0_ROUNDTOINF (
  input      [47:0]   din,
  output     [7:0]    dout
);

  wire       [40:0]   tmp_when_SInt_l131;
  wire       [39:0]   tmp_when_SInt_l137;
  reg        [7:0]    tmp_dout;
  wire                when_SInt_l130;
  wire                when_SInt_l131;
  wire                when_SInt_l137;

  assign tmp_when_SInt_l131 = din[47 : 7];
  assign tmp_when_SInt_l137 = din[46 : 7];
  assign when_SInt_l130 = din[47];
  assign when_SInt_l131 = (! (&tmp_when_SInt_l131));
  always @(*) begin
    if(when_SInt_l130) begin
      if(when_SInt_l131) begin
        tmp_dout = 8'h80;
      end else begin
        tmp_dout = din[7 : 0];
      end
    end else begin
      if(when_SInt_l137) begin
        tmp_dout = 8'h7f;
      end else begin
        tmp_dout = din[7 : 0];
      end
    end
  end

  assign when_SInt_l137 = (|tmp_when_SInt_l137);
  assign dout = tmp_dout;

endmodule

module AMultB (
  input      [29:0]   A,
  input      [17:0]   B,
  output     [47:0]   P,
  input               CEs_0,
  input               CEs_1,
  input               CEs_2,
  input               CEs_3,
  input               clk
);

  wire       [29:0]   dSP48E2_1_ACOUT;
  wire       [17:0]   dSP48E2_1_BCOUT;
  wire       [47:0]   dSP48E2_1_PCOUT;
  wire       [0:0]    dSP48E2_1_CARRYCASCOUT;
  wire       [0:0]    dSP48E2_1_MULTSIGNOUT;
  wire       [47:0]   dSP48E2_1_P;
  wire       [3:0]    dSP48E2_1_CARRYOUT;
  wire       [7:0]    dSP48E2_1_XOROUT;

  DSP48E2 #(
    .A_INPUT("DIRECT"),
    .B_INPUT("DIRECT"),
    .AMULTSEL("A"),
    .BMULTSEL("B"),
    .PREADDINSEL("A"),
    .USE_MULT("MULTIPLY"),
    .USE_SIMD("ONE48"),
    .AREG(2),
    .BREG(2),
    .CREG(1),
    .DREG(1),
    .ADREG(1),
    .MREG(1),
    .PREG(1),
    .ACASCREG(1),
    .BCASCREG(1),
    .CARRYINREG(1),
    .CARRYINSELREG(1),
    .INMODEREG(1),
    .OPMODEREG(1),
    .ALUMODEREG(1) 
  ) dSP48E2_1 (
    .CLK              (clk                      ), //i
    .ALUMODE          (4'b0000                  ), //i
    .INMODE           (5'h0                     ), //i
    .OPMODE           (9'h005                   ), //i
    .CARRYINSEL       (3'b000                   ), //i
    .ACIN             (30'h0                    ), //i
    .BCIN             (18'h0                    ), //i
    .PCIN             (48'h0                    ), //i
    .CARRYCASCIN      (1'b0                     ), //i
    .MULTSIGNIN       (1'b0                     ), //i
    .ACOUT            (dSP48E2_1_ACOUT[29:0]    ), //o
    .BCOUT            (dSP48E2_1_BCOUT[17:0]    ), //o
    .PCOUT            (dSP48E2_1_PCOUT[47:0]    ), //o
    .CARRYCASCOUT     (dSP48E2_1_CARRYCASCOUT   ), //o
    .MULTSIGNOUT      (dSP48E2_1_MULTSIGNOUT    ), //o
    .CEA1             (CEs_0                    ), //i
    .CEA2             (CEs_1                    ), //i
    .CEB1             (CEs_0                    ), //i
    .CEB2             (CEs_1                    ), //i
    .CEC              (1'b0                     ), //i
    .CED              (1'b0                     ), //i
    .CEAD             (1'b0                     ), //i
    .CEM              (CEs_2                    ), //i
    .CEP              (CEs_3                    ), //i
    .CECARRYIN        (1'b0                     ), //i
    .CECTRL           (1'b0                     ), //i
    .CEINMODE         (1'b0                     ), //i
    .CEALUMODE        (1'b0                     ), //i
    .RSTA             (1'b0                     ), //i
    .RSTB             (1'b0                     ), //i
    .RSTC             (1'b0                     ), //i
    .RSTD             (1'b0                     ), //i
    .RSTM             (1'b0                     ), //i
    .RSTP             (1'b0                     ), //i
    .RSTALLCARRYIN    (1'b0                     ), //i
    .RSTCTRL          (1'b0                     ), //i
    .RSTINMODE        (1'b0                     ), //i
    .RSTALUMODE       (1'b0                     ), //i
    .A                (A[29:0]                  ), //i
    .B                (B[17:0]                  ), //i
    .C                (48'h0                    ), //i
    .D                (27'h0                    ), //i
    .CARRYIN          (1'b0                     ), //i
    .P                (dSP48E2_1_P[47:0]        ), //o
    .CARRYOUT         (dSP48E2_1_CARRYOUT[3:0]  ), //o
    .XOROUT           (dSP48E2_1_XOROUT[7:0]    )  //o
  );
  assign P = dSP48E2_1_P;

endmodule

module VideoDownSample (
  input               videoIn_valid,
  output reg          videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 pixCnt;
  reg                 lineCnt;
  wire                pixCntInv;
  wire                lineCntInv;
  wire                fire;
  wire                when_VideoDownSample_l25;
  wire                when_VideoDownSample_l26;
  wire                when_VideoDownSample_l27;
  wire                when_Stream_l408;
  reg                 videoIn_thrown_valid;
  wire                videoIn_thrown_ready;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_0;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_1;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_2;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_3;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_4;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_5;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_6;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_7;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_8;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_9;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_10;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_11;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_12;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_13;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_14;
  wire       [7:0]    videoIn_thrown_payload_frame_line_pixel_15;
  wire                videoIn_thrown_payload_frame_line_endOfLine;
  wire                videoIn_thrown_payload_frame_endOfFrame;
  wire                videoIn_thrown_payload_endOfPack;

  assign pixCntInv = (! pixCnt);
  assign lineCntInv = (! lineCnt);
  assign fire = (videoIn_valid && videoIn_ready);
  assign when_VideoDownSample_l25 = (fire && videoIn_payload_frame_line_endOfLine);
  assign when_VideoDownSample_l26 = (fire && videoIn_payload_frame_line_endOfLine);
  assign when_VideoDownSample_l27 = (fire && videoIn_payload_frame_endOfFrame);
  assign when_Stream_l408 = (pixCnt || lineCnt);
  always @(*) begin
    videoIn_thrown_valid = videoIn_valid;
    if(when_Stream_l408) begin
      videoIn_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    videoIn_ready = videoIn_thrown_ready;
    if(when_Stream_l408) begin
      videoIn_ready = 1'b1;
    end
  end

  assign videoIn_thrown_payload_frame_line_pixel_0 = videoIn_payload_frame_line_pixel_0;
  assign videoIn_thrown_payload_frame_line_pixel_1 = videoIn_payload_frame_line_pixel_1;
  assign videoIn_thrown_payload_frame_line_pixel_2 = videoIn_payload_frame_line_pixel_2;
  assign videoIn_thrown_payload_frame_line_pixel_3 = videoIn_payload_frame_line_pixel_3;
  assign videoIn_thrown_payload_frame_line_pixel_4 = videoIn_payload_frame_line_pixel_4;
  assign videoIn_thrown_payload_frame_line_pixel_5 = videoIn_payload_frame_line_pixel_5;
  assign videoIn_thrown_payload_frame_line_pixel_6 = videoIn_payload_frame_line_pixel_6;
  assign videoIn_thrown_payload_frame_line_pixel_7 = videoIn_payload_frame_line_pixel_7;
  assign videoIn_thrown_payload_frame_line_pixel_8 = videoIn_payload_frame_line_pixel_8;
  assign videoIn_thrown_payload_frame_line_pixel_9 = videoIn_payload_frame_line_pixel_9;
  assign videoIn_thrown_payload_frame_line_pixel_10 = videoIn_payload_frame_line_pixel_10;
  assign videoIn_thrown_payload_frame_line_pixel_11 = videoIn_payload_frame_line_pixel_11;
  assign videoIn_thrown_payload_frame_line_pixel_12 = videoIn_payload_frame_line_pixel_12;
  assign videoIn_thrown_payload_frame_line_pixel_13 = videoIn_payload_frame_line_pixel_13;
  assign videoIn_thrown_payload_frame_line_pixel_14 = videoIn_payload_frame_line_pixel_14;
  assign videoIn_thrown_payload_frame_line_pixel_15 = videoIn_payload_frame_line_pixel_15;
  assign videoIn_thrown_payload_frame_line_endOfLine = videoIn_payload_frame_line_endOfLine;
  assign videoIn_thrown_payload_frame_endOfFrame = videoIn_payload_frame_endOfFrame;
  assign videoIn_thrown_payload_endOfPack = videoIn_payload_endOfPack;
  assign videoOut_valid = videoIn_thrown_valid;
  assign videoIn_thrown_ready = videoOut_ready;
  assign videoOut_payload_frame_line_pixel_0 = videoIn_thrown_payload_frame_line_pixel_0;
  assign videoOut_payload_frame_line_pixel_1 = videoIn_thrown_payload_frame_line_pixel_1;
  assign videoOut_payload_frame_line_pixel_2 = videoIn_thrown_payload_frame_line_pixel_2;
  assign videoOut_payload_frame_line_pixel_3 = videoIn_thrown_payload_frame_line_pixel_3;
  assign videoOut_payload_frame_line_pixel_4 = videoIn_thrown_payload_frame_line_pixel_4;
  assign videoOut_payload_frame_line_pixel_5 = videoIn_thrown_payload_frame_line_pixel_5;
  assign videoOut_payload_frame_line_pixel_6 = videoIn_thrown_payload_frame_line_pixel_6;
  assign videoOut_payload_frame_line_pixel_7 = videoIn_thrown_payload_frame_line_pixel_7;
  assign videoOut_payload_frame_line_pixel_8 = videoIn_thrown_payload_frame_line_pixel_8;
  assign videoOut_payload_frame_line_pixel_9 = videoIn_thrown_payload_frame_line_pixel_9;
  assign videoOut_payload_frame_line_pixel_10 = videoIn_thrown_payload_frame_line_pixel_10;
  assign videoOut_payload_frame_line_pixel_11 = videoIn_thrown_payload_frame_line_pixel_11;
  assign videoOut_payload_frame_line_pixel_12 = videoIn_thrown_payload_frame_line_pixel_12;
  assign videoOut_payload_frame_line_pixel_13 = videoIn_thrown_payload_frame_line_pixel_13;
  assign videoOut_payload_frame_line_pixel_14 = videoIn_thrown_payload_frame_line_pixel_14;
  assign videoOut_payload_frame_line_pixel_15 = videoIn_thrown_payload_frame_line_pixel_15;
  assign videoOut_payload_frame_line_endOfLine = videoIn_thrown_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_endOfFrame = videoIn_thrown_payload_frame_endOfFrame;
  assign videoOut_payload_endOfPack = videoIn_thrown_payload_endOfPack;
  always @(posedge clk) begin
    if(reset) begin
      pixCnt <= 1'b0;
      lineCnt <= 1'b0;
    end else begin
      if(fire) begin
        pixCnt <= pixCntInv;
      end
      if(when_VideoDownSample_l25) begin
        pixCnt <= 1'b0;
      end
      if(when_VideoDownSample_l26) begin
        lineCnt <= lineCntInv;
      end
      if(when_VideoDownSample_l27) begin
        lineCnt <= 1'b0;
      end
    end
  end


endmodule

module SlidingWindowValid (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 line_videoOut_ready;
  reg                 pixel_videoOut_ready;
  wire                line_videoIn_ready;
  wire                line_videoOut_valid;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_0;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_1;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_2;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_3;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_4;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_5;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_6;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_7;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_8;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_9;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_10;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_11;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_12;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_13;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_14;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_0_15;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_0;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_1;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_2;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_3;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_4;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_5;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_6;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_7;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_8;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_9;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_10;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_11;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_12;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_13;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_14;
  wire       [7:0]    line_videoOut_payload_frame_line_pixel_1_15;
  wire                line_videoOut_payload_frame_line_endOfLine;
  wire                line_videoOut_payload_frame_endOfFrame;
  wire                line_videoOut_payload_endOfPack;
  wire                pixel_videoIn_ready;
  wire                pixel_videoOut_valid;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    pixel_videoOut_payload_frame_line_pixel_1_1_15;
  wire                pixel_videoOut_payload_frame_line_endOfLine;
  wire                pixel_videoOut_payload_frame_endOfFrame;
  wire                pixel_videoOut_payload_endOfPack;
  wire                pixelOut_valid;
  wire                pixelOut_ready;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    pixelOut_payload_frame_line_pixel_1_1_15;
  wire                pixelOut_payload_frame_line_endOfLine;
  wire                pixelOut_payload_frame_endOfFrame;
  wire                pixelOut_payload_endOfPack;
  reg                 pixel_videoOut_rValid;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_0_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_0_1_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_0_15;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_0;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_1;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_2;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_3;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_4;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_5;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_6;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_7;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_8;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_9;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_10;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_11;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_12;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_13;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_14;
  reg        [7:0]    pixel_videoOut_rData_frame_line_pixel_1_1_15;
  reg                 pixel_videoOut_rData_frame_line_endOfLine;
  reg                 pixel_videoOut_rData_frame_endOfFrame;
  reg                 pixel_videoOut_rData_endOfPack;
  wire                when_Stream_l342;
  wire                line_videoOut_m2sPipe_valid;
  wire                line_videoOut_m2sPipe_ready;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_0;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_1;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_2;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_3;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_4;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_5;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_6;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_7;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_8;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_9;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_10;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_11;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_12;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_13;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_14;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_0_15;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_0;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_1;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_2;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_3;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_4;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_5;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_6;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_7;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_8;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_9;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_10;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_11;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_12;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_13;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_14;
  wire       [7:0]    line_videoOut_m2sPipe_payload_frame_line_pixel_1_15;
  wire                line_videoOut_m2sPipe_payload_frame_line_endOfLine;
  wire                line_videoOut_m2sPipe_payload_frame_endOfFrame;
  wire                line_videoOut_m2sPipe_payload_endOfPack;
  reg                 line_videoOut_rValid;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_0;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_1;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_2;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_3;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_4;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_5;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_6;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_7;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_8;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_9;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_10;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_11;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_12;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_13;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_14;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_0_15;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_0;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_1;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_2;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_3;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_4;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_5;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_6;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_7;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_8;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_9;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_10;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_11;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_12;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_13;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_14;
  reg        [7:0]    line_videoOut_rData_frame_line_pixel_1_15;
  reg                 line_videoOut_rData_frame_line_endOfLine;
  reg                 line_videoOut_rData_frame_endOfFrame;
  reg                 line_videoOut_rData_endOfPack;
  wire                when_Stream_l342_1;

  LineBufferValid line (
    .videoIn_valid                             (videoIn_valid                                     ), //i
    .videoIn_ready                             (line_videoIn_ready                                ), //o
    .videoIn_payload_frame_line_pixel_0        (videoIn_payload_frame_line_pixel_0[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_1        (videoIn_payload_frame_line_pixel_1[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_2        (videoIn_payload_frame_line_pixel_2[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_3        (videoIn_payload_frame_line_pixel_3[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_4        (videoIn_payload_frame_line_pixel_4[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_5        (videoIn_payload_frame_line_pixel_5[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_6        (videoIn_payload_frame_line_pixel_6[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_7        (videoIn_payload_frame_line_pixel_7[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_8        (videoIn_payload_frame_line_pixel_8[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_9        (videoIn_payload_frame_line_pixel_9[7:0]           ), //i
    .videoIn_payload_frame_line_pixel_10       (videoIn_payload_frame_line_pixel_10[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_11       (videoIn_payload_frame_line_pixel_11[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_12       (videoIn_payload_frame_line_pixel_12[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_13       (videoIn_payload_frame_line_pixel_13[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_14       (videoIn_payload_frame_line_pixel_14[7:0]          ), //i
    .videoIn_payload_frame_line_pixel_15       (videoIn_payload_frame_line_pixel_15[7:0]          ), //i
    .videoIn_payload_frame_line_endOfLine      (videoIn_payload_frame_line_endOfLine              ), //i
    .videoIn_payload_frame_endOfFrame          (videoIn_payload_frame_endOfFrame                  ), //i
    .videoIn_payload_endOfPack                 (videoIn_payload_endOfPack                         ), //i
    .videoOut_valid                            (line_videoOut_valid                               ), //o
    .videoOut_ready                            (line_videoOut_ready                               ), //i
    .videoOut_payload_frame_line_pixel_0_0     (line_videoOut_payload_frame_line_pixel_0_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_1     (line_videoOut_payload_frame_line_pixel_0_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_2     (line_videoOut_payload_frame_line_pixel_0_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_3     (line_videoOut_payload_frame_line_pixel_0_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_4     (line_videoOut_payload_frame_line_pixel_0_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_5     (line_videoOut_payload_frame_line_pixel_0_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_6     (line_videoOut_payload_frame_line_pixel_0_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_7     (line_videoOut_payload_frame_line_pixel_0_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_8     (line_videoOut_payload_frame_line_pixel_0_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_9     (line_videoOut_payload_frame_line_pixel_0_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_0_10    (line_videoOut_payload_frame_line_pixel_0_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_11    (line_videoOut_payload_frame_line_pixel_0_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_12    (line_videoOut_payload_frame_line_pixel_0_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_13    (line_videoOut_payload_frame_line_pixel_0_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_14    (line_videoOut_payload_frame_line_pixel_0_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_0_15    (line_videoOut_payload_frame_line_pixel_0_15[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_0     (line_videoOut_payload_frame_line_pixel_1_0[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_1     (line_videoOut_payload_frame_line_pixel_1_1[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_2     (line_videoOut_payload_frame_line_pixel_1_2[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_3     (line_videoOut_payload_frame_line_pixel_1_3[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_4     (line_videoOut_payload_frame_line_pixel_1_4[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_5     (line_videoOut_payload_frame_line_pixel_1_5[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_6     (line_videoOut_payload_frame_line_pixel_1_6[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_7     (line_videoOut_payload_frame_line_pixel_1_7[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_8     (line_videoOut_payload_frame_line_pixel_1_8[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_9     (line_videoOut_payload_frame_line_pixel_1_9[7:0]   ), //o
    .videoOut_payload_frame_line_pixel_1_10    (line_videoOut_payload_frame_line_pixel_1_10[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_11    (line_videoOut_payload_frame_line_pixel_1_11[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_12    (line_videoOut_payload_frame_line_pixel_1_12[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_13    (line_videoOut_payload_frame_line_pixel_1_13[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_14    (line_videoOut_payload_frame_line_pixel_1_14[7:0]  ), //o
    .videoOut_payload_frame_line_pixel_1_15    (line_videoOut_payload_frame_line_pixel_1_15[7:0]  ), //o
    .videoOut_payload_frame_line_endOfLine     (line_videoOut_payload_frame_line_endOfLine        ), //o
    .videoOut_payload_frame_endOfFrame         (line_videoOut_payload_frame_endOfFrame            ), //o
    .videoOut_payload_endOfPack                (line_videoOut_payload_endOfPack                   ), //o
    .clk                                       (clk                                               ), //i
    .reset                                     (reset                                             )  //i
  );
  PixelBufferValid pixel (
    .videoIn_valid                               (line_videoOut_m2sPipe_valid                               ), //i
    .videoIn_ready                               (pixel_videoIn_ready                                       ), //o
    .videoIn_payload_frame_line_pixel_0_0        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_1        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_2        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_3        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_4        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_5        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_6        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_7        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_8        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_9        (line_videoOut_m2sPipe_payload_frame_line_pixel_0_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_0_10       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_11       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_12       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_13       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_14       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_0_15       (line_videoOut_m2sPipe_payload_frame_line_pixel_0_15[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_0        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_0[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_1        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_1[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_2        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_2[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_3        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_3[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_4        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_4[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_5        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_5[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_6        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_6[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_7        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_7[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_8        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_8[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_9        (line_videoOut_m2sPipe_payload_frame_line_pixel_1_9[7:0]   ), //i
    .videoIn_payload_frame_line_pixel_1_10       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_10[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_11       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_11[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_12       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_12[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_13       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_13[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_14       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_14[7:0]  ), //i
    .videoIn_payload_frame_line_pixel_1_15       (line_videoOut_m2sPipe_payload_frame_line_pixel_1_15[7:0]  ), //i
    .videoIn_payload_frame_line_endOfLine        (line_videoOut_m2sPipe_payload_frame_line_endOfLine        ), //i
    .videoIn_payload_frame_endOfFrame            (line_videoOut_m2sPipe_payload_frame_endOfFrame            ), //i
    .videoIn_payload_endOfPack                   (line_videoOut_m2sPipe_payload_endOfPack                   ), //i
    .videoOut_valid                              (pixel_videoOut_valid                                      ), //o
    .videoOut_ready                              (pixel_videoOut_ready                                      ), //i
    .videoOut_payload_frame_line_pixel_0_0_0     (pixel_videoOut_payload_frame_line_pixel_0_0_0[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_1     (pixel_videoOut_payload_frame_line_pixel_0_0_1[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_2     (pixel_videoOut_payload_frame_line_pixel_0_0_2[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_3     (pixel_videoOut_payload_frame_line_pixel_0_0_3[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_4     (pixel_videoOut_payload_frame_line_pixel_0_0_4[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_5     (pixel_videoOut_payload_frame_line_pixel_0_0_5[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_6     (pixel_videoOut_payload_frame_line_pixel_0_0_6[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_7     (pixel_videoOut_payload_frame_line_pixel_0_0_7[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_8     (pixel_videoOut_payload_frame_line_pixel_0_0_8[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_9     (pixel_videoOut_payload_frame_line_pixel_0_0_9[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_0_10    (pixel_videoOut_payload_frame_line_pixel_0_0_10[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_0_11    (pixel_videoOut_payload_frame_line_pixel_0_0_11[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_0_12    (pixel_videoOut_payload_frame_line_pixel_0_0_12[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_0_13    (pixel_videoOut_payload_frame_line_pixel_0_0_13[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_0_14    (pixel_videoOut_payload_frame_line_pixel_0_0_14[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_0_15    (pixel_videoOut_payload_frame_line_pixel_0_0_15[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_0     (pixel_videoOut_payload_frame_line_pixel_0_1_0[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_1     (pixel_videoOut_payload_frame_line_pixel_0_1_1[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_2     (pixel_videoOut_payload_frame_line_pixel_0_1_2[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_3     (pixel_videoOut_payload_frame_line_pixel_0_1_3[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_4     (pixel_videoOut_payload_frame_line_pixel_0_1_4[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_5     (pixel_videoOut_payload_frame_line_pixel_0_1_5[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_6     (pixel_videoOut_payload_frame_line_pixel_0_1_6[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_7     (pixel_videoOut_payload_frame_line_pixel_0_1_7[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_8     (pixel_videoOut_payload_frame_line_pixel_0_1_8[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_9     (pixel_videoOut_payload_frame_line_pixel_0_1_9[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_0_1_10    (pixel_videoOut_payload_frame_line_pixel_0_1_10[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_11    (pixel_videoOut_payload_frame_line_pixel_0_1_11[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_12    (pixel_videoOut_payload_frame_line_pixel_0_1_12[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_13    (pixel_videoOut_payload_frame_line_pixel_0_1_13[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_14    (pixel_videoOut_payload_frame_line_pixel_0_1_14[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_0_1_15    (pixel_videoOut_payload_frame_line_pixel_0_1_15[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_0     (pixel_videoOut_payload_frame_line_pixel_1_0_0[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_1     (pixel_videoOut_payload_frame_line_pixel_1_0_1[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_2     (pixel_videoOut_payload_frame_line_pixel_1_0_2[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_3     (pixel_videoOut_payload_frame_line_pixel_1_0_3[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_4     (pixel_videoOut_payload_frame_line_pixel_1_0_4[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_5     (pixel_videoOut_payload_frame_line_pixel_1_0_5[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_6     (pixel_videoOut_payload_frame_line_pixel_1_0_6[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_7     (pixel_videoOut_payload_frame_line_pixel_1_0_7[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_8     (pixel_videoOut_payload_frame_line_pixel_1_0_8[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_9     (pixel_videoOut_payload_frame_line_pixel_1_0_9[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_0_10    (pixel_videoOut_payload_frame_line_pixel_1_0_10[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_11    (pixel_videoOut_payload_frame_line_pixel_1_0_11[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_12    (pixel_videoOut_payload_frame_line_pixel_1_0_12[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_13    (pixel_videoOut_payload_frame_line_pixel_1_0_13[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_14    (pixel_videoOut_payload_frame_line_pixel_1_0_14[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_0_15    (pixel_videoOut_payload_frame_line_pixel_1_0_15[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_0     (pixel_videoOut_payload_frame_line_pixel_1_1_0[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_1     (pixel_videoOut_payload_frame_line_pixel_1_1_1[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_2     (pixel_videoOut_payload_frame_line_pixel_1_1_2[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_3     (pixel_videoOut_payload_frame_line_pixel_1_1_3[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_4     (pixel_videoOut_payload_frame_line_pixel_1_1_4[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_5     (pixel_videoOut_payload_frame_line_pixel_1_1_5[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_6     (pixel_videoOut_payload_frame_line_pixel_1_1_6[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_7     (pixel_videoOut_payload_frame_line_pixel_1_1_7[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_8     (pixel_videoOut_payload_frame_line_pixel_1_1_8[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_9     (pixel_videoOut_payload_frame_line_pixel_1_1_9[7:0]        ), //o
    .videoOut_payload_frame_line_pixel_1_1_10    (pixel_videoOut_payload_frame_line_pixel_1_1_10[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_11    (pixel_videoOut_payload_frame_line_pixel_1_1_11[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_12    (pixel_videoOut_payload_frame_line_pixel_1_1_12[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_13    (pixel_videoOut_payload_frame_line_pixel_1_1_13[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_14    (pixel_videoOut_payload_frame_line_pixel_1_1_14[7:0]       ), //o
    .videoOut_payload_frame_line_pixel_1_1_15    (pixel_videoOut_payload_frame_line_pixel_1_1_15[7:0]       ), //o
    .videoOut_payload_frame_line_endOfLine       (pixel_videoOut_payload_frame_line_endOfLine               ), //o
    .videoOut_payload_frame_endOfFrame           (pixel_videoOut_payload_frame_endOfFrame                   ), //o
    .videoOut_payload_endOfPack                  (pixel_videoOut_payload_endOfPack                          ), //o
    .clk                                         (clk                                                       ), //i
    .reset                                       (reset                                                     )  //i
  );
  always @(*) begin
    pixel_videoOut_ready = pixelOut_ready;
    if(when_Stream_l342) begin
      pixel_videoOut_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! pixelOut_valid);
  assign pixelOut_valid = pixel_videoOut_rValid;
  assign pixelOut_payload_frame_line_pixel_0_0_0 = pixel_videoOut_rData_frame_line_pixel_0_0_0;
  assign pixelOut_payload_frame_line_pixel_0_0_1 = pixel_videoOut_rData_frame_line_pixel_0_0_1;
  assign pixelOut_payload_frame_line_pixel_0_0_2 = pixel_videoOut_rData_frame_line_pixel_0_0_2;
  assign pixelOut_payload_frame_line_pixel_0_0_3 = pixel_videoOut_rData_frame_line_pixel_0_0_3;
  assign pixelOut_payload_frame_line_pixel_0_0_4 = pixel_videoOut_rData_frame_line_pixel_0_0_4;
  assign pixelOut_payload_frame_line_pixel_0_0_5 = pixel_videoOut_rData_frame_line_pixel_0_0_5;
  assign pixelOut_payload_frame_line_pixel_0_0_6 = pixel_videoOut_rData_frame_line_pixel_0_0_6;
  assign pixelOut_payload_frame_line_pixel_0_0_7 = pixel_videoOut_rData_frame_line_pixel_0_0_7;
  assign pixelOut_payload_frame_line_pixel_0_0_8 = pixel_videoOut_rData_frame_line_pixel_0_0_8;
  assign pixelOut_payload_frame_line_pixel_0_0_9 = pixel_videoOut_rData_frame_line_pixel_0_0_9;
  assign pixelOut_payload_frame_line_pixel_0_0_10 = pixel_videoOut_rData_frame_line_pixel_0_0_10;
  assign pixelOut_payload_frame_line_pixel_0_0_11 = pixel_videoOut_rData_frame_line_pixel_0_0_11;
  assign pixelOut_payload_frame_line_pixel_0_0_12 = pixel_videoOut_rData_frame_line_pixel_0_0_12;
  assign pixelOut_payload_frame_line_pixel_0_0_13 = pixel_videoOut_rData_frame_line_pixel_0_0_13;
  assign pixelOut_payload_frame_line_pixel_0_0_14 = pixel_videoOut_rData_frame_line_pixel_0_0_14;
  assign pixelOut_payload_frame_line_pixel_0_0_15 = pixel_videoOut_rData_frame_line_pixel_0_0_15;
  assign pixelOut_payload_frame_line_pixel_0_1_0 = pixel_videoOut_rData_frame_line_pixel_0_1_0;
  assign pixelOut_payload_frame_line_pixel_0_1_1 = pixel_videoOut_rData_frame_line_pixel_0_1_1;
  assign pixelOut_payload_frame_line_pixel_0_1_2 = pixel_videoOut_rData_frame_line_pixel_0_1_2;
  assign pixelOut_payload_frame_line_pixel_0_1_3 = pixel_videoOut_rData_frame_line_pixel_0_1_3;
  assign pixelOut_payload_frame_line_pixel_0_1_4 = pixel_videoOut_rData_frame_line_pixel_0_1_4;
  assign pixelOut_payload_frame_line_pixel_0_1_5 = pixel_videoOut_rData_frame_line_pixel_0_1_5;
  assign pixelOut_payload_frame_line_pixel_0_1_6 = pixel_videoOut_rData_frame_line_pixel_0_1_6;
  assign pixelOut_payload_frame_line_pixel_0_1_7 = pixel_videoOut_rData_frame_line_pixel_0_1_7;
  assign pixelOut_payload_frame_line_pixel_0_1_8 = pixel_videoOut_rData_frame_line_pixel_0_1_8;
  assign pixelOut_payload_frame_line_pixel_0_1_9 = pixel_videoOut_rData_frame_line_pixel_0_1_9;
  assign pixelOut_payload_frame_line_pixel_0_1_10 = pixel_videoOut_rData_frame_line_pixel_0_1_10;
  assign pixelOut_payload_frame_line_pixel_0_1_11 = pixel_videoOut_rData_frame_line_pixel_0_1_11;
  assign pixelOut_payload_frame_line_pixel_0_1_12 = pixel_videoOut_rData_frame_line_pixel_0_1_12;
  assign pixelOut_payload_frame_line_pixel_0_1_13 = pixel_videoOut_rData_frame_line_pixel_0_1_13;
  assign pixelOut_payload_frame_line_pixel_0_1_14 = pixel_videoOut_rData_frame_line_pixel_0_1_14;
  assign pixelOut_payload_frame_line_pixel_0_1_15 = pixel_videoOut_rData_frame_line_pixel_0_1_15;
  assign pixelOut_payload_frame_line_pixel_1_0_0 = pixel_videoOut_rData_frame_line_pixel_1_0_0;
  assign pixelOut_payload_frame_line_pixel_1_0_1 = pixel_videoOut_rData_frame_line_pixel_1_0_1;
  assign pixelOut_payload_frame_line_pixel_1_0_2 = pixel_videoOut_rData_frame_line_pixel_1_0_2;
  assign pixelOut_payload_frame_line_pixel_1_0_3 = pixel_videoOut_rData_frame_line_pixel_1_0_3;
  assign pixelOut_payload_frame_line_pixel_1_0_4 = pixel_videoOut_rData_frame_line_pixel_1_0_4;
  assign pixelOut_payload_frame_line_pixel_1_0_5 = pixel_videoOut_rData_frame_line_pixel_1_0_5;
  assign pixelOut_payload_frame_line_pixel_1_0_6 = pixel_videoOut_rData_frame_line_pixel_1_0_6;
  assign pixelOut_payload_frame_line_pixel_1_0_7 = pixel_videoOut_rData_frame_line_pixel_1_0_7;
  assign pixelOut_payload_frame_line_pixel_1_0_8 = pixel_videoOut_rData_frame_line_pixel_1_0_8;
  assign pixelOut_payload_frame_line_pixel_1_0_9 = pixel_videoOut_rData_frame_line_pixel_1_0_9;
  assign pixelOut_payload_frame_line_pixel_1_0_10 = pixel_videoOut_rData_frame_line_pixel_1_0_10;
  assign pixelOut_payload_frame_line_pixel_1_0_11 = pixel_videoOut_rData_frame_line_pixel_1_0_11;
  assign pixelOut_payload_frame_line_pixel_1_0_12 = pixel_videoOut_rData_frame_line_pixel_1_0_12;
  assign pixelOut_payload_frame_line_pixel_1_0_13 = pixel_videoOut_rData_frame_line_pixel_1_0_13;
  assign pixelOut_payload_frame_line_pixel_1_0_14 = pixel_videoOut_rData_frame_line_pixel_1_0_14;
  assign pixelOut_payload_frame_line_pixel_1_0_15 = pixel_videoOut_rData_frame_line_pixel_1_0_15;
  assign pixelOut_payload_frame_line_pixel_1_1_0 = pixel_videoOut_rData_frame_line_pixel_1_1_0;
  assign pixelOut_payload_frame_line_pixel_1_1_1 = pixel_videoOut_rData_frame_line_pixel_1_1_1;
  assign pixelOut_payload_frame_line_pixel_1_1_2 = pixel_videoOut_rData_frame_line_pixel_1_1_2;
  assign pixelOut_payload_frame_line_pixel_1_1_3 = pixel_videoOut_rData_frame_line_pixel_1_1_3;
  assign pixelOut_payload_frame_line_pixel_1_1_4 = pixel_videoOut_rData_frame_line_pixel_1_1_4;
  assign pixelOut_payload_frame_line_pixel_1_1_5 = pixel_videoOut_rData_frame_line_pixel_1_1_5;
  assign pixelOut_payload_frame_line_pixel_1_1_6 = pixel_videoOut_rData_frame_line_pixel_1_1_6;
  assign pixelOut_payload_frame_line_pixel_1_1_7 = pixel_videoOut_rData_frame_line_pixel_1_1_7;
  assign pixelOut_payload_frame_line_pixel_1_1_8 = pixel_videoOut_rData_frame_line_pixel_1_1_8;
  assign pixelOut_payload_frame_line_pixel_1_1_9 = pixel_videoOut_rData_frame_line_pixel_1_1_9;
  assign pixelOut_payload_frame_line_pixel_1_1_10 = pixel_videoOut_rData_frame_line_pixel_1_1_10;
  assign pixelOut_payload_frame_line_pixel_1_1_11 = pixel_videoOut_rData_frame_line_pixel_1_1_11;
  assign pixelOut_payload_frame_line_pixel_1_1_12 = pixel_videoOut_rData_frame_line_pixel_1_1_12;
  assign pixelOut_payload_frame_line_pixel_1_1_13 = pixel_videoOut_rData_frame_line_pixel_1_1_13;
  assign pixelOut_payload_frame_line_pixel_1_1_14 = pixel_videoOut_rData_frame_line_pixel_1_1_14;
  assign pixelOut_payload_frame_line_pixel_1_1_15 = pixel_videoOut_rData_frame_line_pixel_1_1_15;
  assign pixelOut_payload_frame_line_endOfLine = pixel_videoOut_rData_frame_line_endOfLine;
  assign pixelOut_payload_frame_endOfFrame = pixel_videoOut_rData_frame_endOfFrame;
  assign pixelOut_payload_endOfPack = pixel_videoOut_rData_endOfPack;
  assign videoIn_ready = line_videoIn_ready;
  always @(*) begin
    line_videoOut_ready = line_videoOut_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      line_videoOut_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! line_videoOut_m2sPipe_valid);
  assign line_videoOut_m2sPipe_valid = line_videoOut_rValid;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_0 = line_videoOut_rData_frame_line_pixel_0_0;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_1 = line_videoOut_rData_frame_line_pixel_0_1;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_2 = line_videoOut_rData_frame_line_pixel_0_2;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_3 = line_videoOut_rData_frame_line_pixel_0_3;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_4 = line_videoOut_rData_frame_line_pixel_0_4;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_5 = line_videoOut_rData_frame_line_pixel_0_5;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_6 = line_videoOut_rData_frame_line_pixel_0_6;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_7 = line_videoOut_rData_frame_line_pixel_0_7;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_8 = line_videoOut_rData_frame_line_pixel_0_8;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_9 = line_videoOut_rData_frame_line_pixel_0_9;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_10 = line_videoOut_rData_frame_line_pixel_0_10;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_11 = line_videoOut_rData_frame_line_pixel_0_11;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_12 = line_videoOut_rData_frame_line_pixel_0_12;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_13 = line_videoOut_rData_frame_line_pixel_0_13;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_14 = line_videoOut_rData_frame_line_pixel_0_14;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_0_15 = line_videoOut_rData_frame_line_pixel_0_15;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_0 = line_videoOut_rData_frame_line_pixel_1_0;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_1 = line_videoOut_rData_frame_line_pixel_1_1;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_2 = line_videoOut_rData_frame_line_pixel_1_2;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_3 = line_videoOut_rData_frame_line_pixel_1_3;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_4 = line_videoOut_rData_frame_line_pixel_1_4;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_5 = line_videoOut_rData_frame_line_pixel_1_5;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_6 = line_videoOut_rData_frame_line_pixel_1_6;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_7 = line_videoOut_rData_frame_line_pixel_1_7;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_8 = line_videoOut_rData_frame_line_pixel_1_8;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_9 = line_videoOut_rData_frame_line_pixel_1_9;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_10 = line_videoOut_rData_frame_line_pixel_1_10;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_11 = line_videoOut_rData_frame_line_pixel_1_11;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_12 = line_videoOut_rData_frame_line_pixel_1_12;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_13 = line_videoOut_rData_frame_line_pixel_1_13;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_14 = line_videoOut_rData_frame_line_pixel_1_14;
  assign line_videoOut_m2sPipe_payload_frame_line_pixel_1_15 = line_videoOut_rData_frame_line_pixel_1_15;
  assign line_videoOut_m2sPipe_payload_frame_line_endOfLine = line_videoOut_rData_frame_line_endOfLine;
  assign line_videoOut_m2sPipe_payload_frame_endOfFrame = line_videoOut_rData_frame_endOfFrame;
  assign line_videoOut_m2sPipe_payload_endOfPack = line_videoOut_rData_endOfPack;
  assign line_videoOut_m2sPipe_ready = pixel_videoIn_ready;
  assign videoOut_valid = pixelOut_valid;
  assign pixelOut_ready = videoOut_ready;
  assign videoOut_payload_endOfPack = pixelOut_payload_endOfPack;
  assign videoOut_payload_frame_endOfFrame = pixelOut_payload_frame_endOfFrame;
  assign videoOut_payload_frame_line_endOfLine = pixelOut_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_line_pixel_0_0_0 = pixelOut_payload_frame_line_pixel_0_0_0;
  assign videoOut_payload_frame_line_pixel_0_0_1 = pixelOut_payload_frame_line_pixel_0_0_1;
  assign videoOut_payload_frame_line_pixel_0_0_2 = pixelOut_payload_frame_line_pixel_0_0_2;
  assign videoOut_payload_frame_line_pixel_0_0_3 = pixelOut_payload_frame_line_pixel_0_0_3;
  assign videoOut_payload_frame_line_pixel_0_0_4 = pixelOut_payload_frame_line_pixel_0_0_4;
  assign videoOut_payload_frame_line_pixel_0_0_5 = pixelOut_payload_frame_line_pixel_0_0_5;
  assign videoOut_payload_frame_line_pixel_0_0_6 = pixelOut_payload_frame_line_pixel_0_0_6;
  assign videoOut_payload_frame_line_pixel_0_0_7 = pixelOut_payload_frame_line_pixel_0_0_7;
  assign videoOut_payload_frame_line_pixel_0_0_8 = pixelOut_payload_frame_line_pixel_0_0_8;
  assign videoOut_payload_frame_line_pixel_0_0_9 = pixelOut_payload_frame_line_pixel_0_0_9;
  assign videoOut_payload_frame_line_pixel_0_0_10 = pixelOut_payload_frame_line_pixel_0_0_10;
  assign videoOut_payload_frame_line_pixel_0_0_11 = pixelOut_payload_frame_line_pixel_0_0_11;
  assign videoOut_payload_frame_line_pixel_0_0_12 = pixelOut_payload_frame_line_pixel_0_0_12;
  assign videoOut_payload_frame_line_pixel_0_0_13 = pixelOut_payload_frame_line_pixel_0_0_13;
  assign videoOut_payload_frame_line_pixel_0_0_14 = pixelOut_payload_frame_line_pixel_0_0_14;
  assign videoOut_payload_frame_line_pixel_0_0_15 = pixelOut_payload_frame_line_pixel_0_0_15;
  assign videoOut_payload_frame_line_pixel_0_1_0 = pixelOut_payload_frame_line_pixel_1_0_0;
  assign videoOut_payload_frame_line_pixel_0_1_1 = pixelOut_payload_frame_line_pixel_1_0_1;
  assign videoOut_payload_frame_line_pixel_0_1_2 = pixelOut_payload_frame_line_pixel_1_0_2;
  assign videoOut_payload_frame_line_pixel_0_1_3 = pixelOut_payload_frame_line_pixel_1_0_3;
  assign videoOut_payload_frame_line_pixel_0_1_4 = pixelOut_payload_frame_line_pixel_1_0_4;
  assign videoOut_payload_frame_line_pixel_0_1_5 = pixelOut_payload_frame_line_pixel_1_0_5;
  assign videoOut_payload_frame_line_pixel_0_1_6 = pixelOut_payload_frame_line_pixel_1_0_6;
  assign videoOut_payload_frame_line_pixel_0_1_7 = pixelOut_payload_frame_line_pixel_1_0_7;
  assign videoOut_payload_frame_line_pixel_0_1_8 = pixelOut_payload_frame_line_pixel_1_0_8;
  assign videoOut_payload_frame_line_pixel_0_1_9 = pixelOut_payload_frame_line_pixel_1_0_9;
  assign videoOut_payload_frame_line_pixel_0_1_10 = pixelOut_payload_frame_line_pixel_1_0_10;
  assign videoOut_payload_frame_line_pixel_0_1_11 = pixelOut_payload_frame_line_pixel_1_0_11;
  assign videoOut_payload_frame_line_pixel_0_1_12 = pixelOut_payload_frame_line_pixel_1_0_12;
  assign videoOut_payload_frame_line_pixel_0_1_13 = pixelOut_payload_frame_line_pixel_1_0_13;
  assign videoOut_payload_frame_line_pixel_0_1_14 = pixelOut_payload_frame_line_pixel_1_0_14;
  assign videoOut_payload_frame_line_pixel_0_1_15 = pixelOut_payload_frame_line_pixel_1_0_15;
  assign videoOut_payload_frame_line_pixel_1_0_0 = pixelOut_payload_frame_line_pixel_0_1_0;
  assign videoOut_payload_frame_line_pixel_1_0_1 = pixelOut_payload_frame_line_pixel_0_1_1;
  assign videoOut_payload_frame_line_pixel_1_0_2 = pixelOut_payload_frame_line_pixel_0_1_2;
  assign videoOut_payload_frame_line_pixel_1_0_3 = pixelOut_payload_frame_line_pixel_0_1_3;
  assign videoOut_payload_frame_line_pixel_1_0_4 = pixelOut_payload_frame_line_pixel_0_1_4;
  assign videoOut_payload_frame_line_pixel_1_0_5 = pixelOut_payload_frame_line_pixel_0_1_5;
  assign videoOut_payload_frame_line_pixel_1_0_6 = pixelOut_payload_frame_line_pixel_0_1_6;
  assign videoOut_payload_frame_line_pixel_1_0_7 = pixelOut_payload_frame_line_pixel_0_1_7;
  assign videoOut_payload_frame_line_pixel_1_0_8 = pixelOut_payload_frame_line_pixel_0_1_8;
  assign videoOut_payload_frame_line_pixel_1_0_9 = pixelOut_payload_frame_line_pixel_0_1_9;
  assign videoOut_payload_frame_line_pixel_1_0_10 = pixelOut_payload_frame_line_pixel_0_1_10;
  assign videoOut_payload_frame_line_pixel_1_0_11 = pixelOut_payload_frame_line_pixel_0_1_11;
  assign videoOut_payload_frame_line_pixel_1_0_12 = pixelOut_payload_frame_line_pixel_0_1_12;
  assign videoOut_payload_frame_line_pixel_1_0_13 = pixelOut_payload_frame_line_pixel_0_1_13;
  assign videoOut_payload_frame_line_pixel_1_0_14 = pixelOut_payload_frame_line_pixel_0_1_14;
  assign videoOut_payload_frame_line_pixel_1_0_15 = pixelOut_payload_frame_line_pixel_0_1_15;
  assign videoOut_payload_frame_line_pixel_1_1_0 = pixelOut_payload_frame_line_pixel_1_1_0;
  assign videoOut_payload_frame_line_pixel_1_1_1 = pixelOut_payload_frame_line_pixel_1_1_1;
  assign videoOut_payload_frame_line_pixel_1_1_2 = pixelOut_payload_frame_line_pixel_1_1_2;
  assign videoOut_payload_frame_line_pixel_1_1_3 = pixelOut_payload_frame_line_pixel_1_1_3;
  assign videoOut_payload_frame_line_pixel_1_1_4 = pixelOut_payload_frame_line_pixel_1_1_4;
  assign videoOut_payload_frame_line_pixel_1_1_5 = pixelOut_payload_frame_line_pixel_1_1_5;
  assign videoOut_payload_frame_line_pixel_1_1_6 = pixelOut_payload_frame_line_pixel_1_1_6;
  assign videoOut_payload_frame_line_pixel_1_1_7 = pixelOut_payload_frame_line_pixel_1_1_7;
  assign videoOut_payload_frame_line_pixel_1_1_8 = pixelOut_payload_frame_line_pixel_1_1_8;
  assign videoOut_payload_frame_line_pixel_1_1_9 = pixelOut_payload_frame_line_pixel_1_1_9;
  assign videoOut_payload_frame_line_pixel_1_1_10 = pixelOut_payload_frame_line_pixel_1_1_10;
  assign videoOut_payload_frame_line_pixel_1_1_11 = pixelOut_payload_frame_line_pixel_1_1_11;
  assign videoOut_payload_frame_line_pixel_1_1_12 = pixelOut_payload_frame_line_pixel_1_1_12;
  assign videoOut_payload_frame_line_pixel_1_1_13 = pixelOut_payload_frame_line_pixel_1_1_13;
  assign videoOut_payload_frame_line_pixel_1_1_14 = pixelOut_payload_frame_line_pixel_1_1_14;
  assign videoOut_payload_frame_line_pixel_1_1_15 = pixelOut_payload_frame_line_pixel_1_1_15;
  always @(posedge clk) begin
    if(reset) begin
      pixel_videoOut_rValid <= 1'b0;
      line_videoOut_rValid <= 1'b0;
    end else begin
      if(pixel_videoOut_ready) begin
        pixel_videoOut_rValid <= pixel_videoOut_valid;
      end
      if(line_videoOut_ready) begin
        line_videoOut_rValid <= line_videoOut_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(pixel_videoOut_ready) begin
      pixel_videoOut_rData_frame_line_pixel_0_0_0 <= pixel_videoOut_payload_frame_line_pixel_0_0_0;
      pixel_videoOut_rData_frame_line_pixel_0_0_1 <= pixel_videoOut_payload_frame_line_pixel_0_0_1;
      pixel_videoOut_rData_frame_line_pixel_0_0_2 <= pixel_videoOut_payload_frame_line_pixel_0_0_2;
      pixel_videoOut_rData_frame_line_pixel_0_0_3 <= pixel_videoOut_payload_frame_line_pixel_0_0_3;
      pixel_videoOut_rData_frame_line_pixel_0_0_4 <= pixel_videoOut_payload_frame_line_pixel_0_0_4;
      pixel_videoOut_rData_frame_line_pixel_0_0_5 <= pixel_videoOut_payload_frame_line_pixel_0_0_5;
      pixel_videoOut_rData_frame_line_pixel_0_0_6 <= pixel_videoOut_payload_frame_line_pixel_0_0_6;
      pixel_videoOut_rData_frame_line_pixel_0_0_7 <= pixel_videoOut_payload_frame_line_pixel_0_0_7;
      pixel_videoOut_rData_frame_line_pixel_0_0_8 <= pixel_videoOut_payload_frame_line_pixel_0_0_8;
      pixel_videoOut_rData_frame_line_pixel_0_0_9 <= pixel_videoOut_payload_frame_line_pixel_0_0_9;
      pixel_videoOut_rData_frame_line_pixel_0_0_10 <= pixel_videoOut_payload_frame_line_pixel_0_0_10;
      pixel_videoOut_rData_frame_line_pixel_0_0_11 <= pixel_videoOut_payload_frame_line_pixel_0_0_11;
      pixel_videoOut_rData_frame_line_pixel_0_0_12 <= pixel_videoOut_payload_frame_line_pixel_0_0_12;
      pixel_videoOut_rData_frame_line_pixel_0_0_13 <= pixel_videoOut_payload_frame_line_pixel_0_0_13;
      pixel_videoOut_rData_frame_line_pixel_0_0_14 <= pixel_videoOut_payload_frame_line_pixel_0_0_14;
      pixel_videoOut_rData_frame_line_pixel_0_0_15 <= pixel_videoOut_payload_frame_line_pixel_0_0_15;
      pixel_videoOut_rData_frame_line_pixel_0_1_0 <= pixel_videoOut_payload_frame_line_pixel_0_1_0;
      pixel_videoOut_rData_frame_line_pixel_0_1_1 <= pixel_videoOut_payload_frame_line_pixel_0_1_1;
      pixel_videoOut_rData_frame_line_pixel_0_1_2 <= pixel_videoOut_payload_frame_line_pixel_0_1_2;
      pixel_videoOut_rData_frame_line_pixel_0_1_3 <= pixel_videoOut_payload_frame_line_pixel_0_1_3;
      pixel_videoOut_rData_frame_line_pixel_0_1_4 <= pixel_videoOut_payload_frame_line_pixel_0_1_4;
      pixel_videoOut_rData_frame_line_pixel_0_1_5 <= pixel_videoOut_payload_frame_line_pixel_0_1_5;
      pixel_videoOut_rData_frame_line_pixel_0_1_6 <= pixel_videoOut_payload_frame_line_pixel_0_1_6;
      pixel_videoOut_rData_frame_line_pixel_0_1_7 <= pixel_videoOut_payload_frame_line_pixel_0_1_7;
      pixel_videoOut_rData_frame_line_pixel_0_1_8 <= pixel_videoOut_payload_frame_line_pixel_0_1_8;
      pixel_videoOut_rData_frame_line_pixel_0_1_9 <= pixel_videoOut_payload_frame_line_pixel_0_1_9;
      pixel_videoOut_rData_frame_line_pixel_0_1_10 <= pixel_videoOut_payload_frame_line_pixel_0_1_10;
      pixel_videoOut_rData_frame_line_pixel_0_1_11 <= pixel_videoOut_payload_frame_line_pixel_0_1_11;
      pixel_videoOut_rData_frame_line_pixel_0_1_12 <= pixel_videoOut_payload_frame_line_pixel_0_1_12;
      pixel_videoOut_rData_frame_line_pixel_0_1_13 <= pixel_videoOut_payload_frame_line_pixel_0_1_13;
      pixel_videoOut_rData_frame_line_pixel_0_1_14 <= pixel_videoOut_payload_frame_line_pixel_0_1_14;
      pixel_videoOut_rData_frame_line_pixel_0_1_15 <= pixel_videoOut_payload_frame_line_pixel_0_1_15;
      pixel_videoOut_rData_frame_line_pixel_1_0_0 <= pixel_videoOut_payload_frame_line_pixel_1_0_0;
      pixel_videoOut_rData_frame_line_pixel_1_0_1 <= pixel_videoOut_payload_frame_line_pixel_1_0_1;
      pixel_videoOut_rData_frame_line_pixel_1_0_2 <= pixel_videoOut_payload_frame_line_pixel_1_0_2;
      pixel_videoOut_rData_frame_line_pixel_1_0_3 <= pixel_videoOut_payload_frame_line_pixel_1_0_3;
      pixel_videoOut_rData_frame_line_pixel_1_0_4 <= pixel_videoOut_payload_frame_line_pixel_1_0_4;
      pixel_videoOut_rData_frame_line_pixel_1_0_5 <= pixel_videoOut_payload_frame_line_pixel_1_0_5;
      pixel_videoOut_rData_frame_line_pixel_1_0_6 <= pixel_videoOut_payload_frame_line_pixel_1_0_6;
      pixel_videoOut_rData_frame_line_pixel_1_0_7 <= pixel_videoOut_payload_frame_line_pixel_1_0_7;
      pixel_videoOut_rData_frame_line_pixel_1_0_8 <= pixel_videoOut_payload_frame_line_pixel_1_0_8;
      pixel_videoOut_rData_frame_line_pixel_1_0_9 <= pixel_videoOut_payload_frame_line_pixel_1_0_9;
      pixel_videoOut_rData_frame_line_pixel_1_0_10 <= pixel_videoOut_payload_frame_line_pixel_1_0_10;
      pixel_videoOut_rData_frame_line_pixel_1_0_11 <= pixel_videoOut_payload_frame_line_pixel_1_0_11;
      pixel_videoOut_rData_frame_line_pixel_1_0_12 <= pixel_videoOut_payload_frame_line_pixel_1_0_12;
      pixel_videoOut_rData_frame_line_pixel_1_0_13 <= pixel_videoOut_payload_frame_line_pixel_1_0_13;
      pixel_videoOut_rData_frame_line_pixel_1_0_14 <= pixel_videoOut_payload_frame_line_pixel_1_0_14;
      pixel_videoOut_rData_frame_line_pixel_1_0_15 <= pixel_videoOut_payload_frame_line_pixel_1_0_15;
      pixel_videoOut_rData_frame_line_pixel_1_1_0 <= pixel_videoOut_payload_frame_line_pixel_1_1_0;
      pixel_videoOut_rData_frame_line_pixel_1_1_1 <= pixel_videoOut_payload_frame_line_pixel_1_1_1;
      pixel_videoOut_rData_frame_line_pixel_1_1_2 <= pixel_videoOut_payload_frame_line_pixel_1_1_2;
      pixel_videoOut_rData_frame_line_pixel_1_1_3 <= pixel_videoOut_payload_frame_line_pixel_1_1_3;
      pixel_videoOut_rData_frame_line_pixel_1_1_4 <= pixel_videoOut_payload_frame_line_pixel_1_1_4;
      pixel_videoOut_rData_frame_line_pixel_1_1_5 <= pixel_videoOut_payload_frame_line_pixel_1_1_5;
      pixel_videoOut_rData_frame_line_pixel_1_1_6 <= pixel_videoOut_payload_frame_line_pixel_1_1_6;
      pixel_videoOut_rData_frame_line_pixel_1_1_7 <= pixel_videoOut_payload_frame_line_pixel_1_1_7;
      pixel_videoOut_rData_frame_line_pixel_1_1_8 <= pixel_videoOut_payload_frame_line_pixel_1_1_8;
      pixel_videoOut_rData_frame_line_pixel_1_1_9 <= pixel_videoOut_payload_frame_line_pixel_1_1_9;
      pixel_videoOut_rData_frame_line_pixel_1_1_10 <= pixel_videoOut_payload_frame_line_pixel_1_1_10;
      pixel_videoOut_rData_frame_line_pixel_1_1_11 <= pixel_videoOut_payload_frame_line_pixel_1_1_11;
      pixel_videoOut_rData_frame_line_pixel_1_1_12 <= pixel_videoOut_payload_frame_line_pixel_1_1_12;
      pixel_videoOut_rData_frame_line_pixel_1_1_13 <= pixel_videoOut_payload_frame_line_pixel_1_1_13;
      pixel_videoOut_rData_frame_line_pixel_1_1_14 <= pixel_videoOut_payload_frame_line_pixel_1_1_14;
      pixel_videoOut_rData_frame_line_pixel_1_1_15 <= pixel_videoOut_payload_frame_line_pixel_1_1_15;
      pixel_videoOut_rData_frame_line_endOfLine <= pixel_videoOut_payload_frame_line_endOfLine;
      pixel_videoOut_rData_frame_endOfFrame <= pixel_videoOut_payload_frame_endOfFrame;
      pixel_videoOut_rData_endOfPack <= pixel_videoOut_payload_endOfPack;
    end
    if(line_videoOut_ready) begin
      line_videoOut_rData_frame_line_pixel_0_0 <= line_videoOut_payload_frame_line_pixel_0_0;
      line_videoOut_rData_frame_line_pixel_0_1 <= line_videoOut_payload_frame_line_pixel_0_1;
      line_videoOut_rData_frame_line_pixel_0_2 <= line_videoOut_payload_frame_line_pixel_0_2;
      line_videoOut_rData_frame_line_pixel_0_3 <= line_videoOut_payload_frame_line_pixel_0_3;
      line_videoOut_rData_frame_line_pixel_0_4 <= line_videoOut_payload_frame_line_pixel_0_4;
      line_videoOut_rData_frame_line_pixel_0_5 <= line_videoOut_payload_frame_line_pixel_0_5;
      line_videoOut_rData_frame_line_pixel_0_6 <= line_videoOut_payload_frame_line_pixel_0_6;
      line_videoOut_rData_frame_line_pixel_0_7 <= line_videoOut_payload_frame_line_pixel_0_7;
      line_videoOut_rData_frame_line_pixel_0_8 <= line_videoOut_payload_frame_line_pixel_0_8;
      line_videoOut_rData_frame_line_pixel_0_9 <= line_videoOut_payload_frame_line_pixel_0_9;
      line_videoOut_rData_frame_line_pixel_0_10 <= line_videoOut_payload_frame_line_pixel_0_10;
      line_videoOut_rData_frame_line_pixel_0_11 <= line_videoOut_payload_frame_line_pixel_0_11;
      line_videoOut_rData_frame_line_pixel_0_12 <= line_videoOut_payload_frame_line_pixel_0_12;
      line_videoOut_rData_frame_line_pixel_0_13 <= line_videoOut_payload_frame_line_pixel_0_13;
      line_videoOut_rData_frame_line_pixel_0_14 <= line_videoOut_payload_frame_line_pixel_0_14;
      line_videoOut_rData_frame_line_pixel_0_15 <= line_videoOut_payload_frame_line_pixel_0_15;
      line_videoOut_rData_frame_line_pixel_1_0 <= line_videoOut_payload_frame_line_pixel_1_0;
      line_videoOut_rData_frame_line_pixel_1_1 <= line_videoOut_payload_frame_line_pixel_1_1;
      line_videoOut_rData_frame_line_pixel_1_2 <= line_videoOut_payload_frame_line_pixel_1_2;
      line_videoOut_rData_frame_line_pixel_1_3 <= line_videoOut_payload_frame_line_pixel_1_3;
      line_videoOut_rData_frame_line_pixel_1_4 <= line_videoOut_payload_frame_line_pixel_1_4;
      line_videoOut_rData_frame_line_pixel_1_5 <= line_videoOut_payload_frame_line_pixel_1_5;
      line_videoOut_rData_frame_line_pixel_1_6 <= line_videoOut_payload_frame_line_pixel_1_6;
      line_videoOut_rData_frame_line_pixel_1_7 <= line_videoOut_payload_frame_line_pixel_1_7;
      line_videoOut_rData_frame_line_pixel_1_8 <= line_videoOut_payload_frame_line_pixel_1_8;
      line_videoOut_rData_frame_line_pixel_1_9 <= line_videoOut_payload_frame_line_pixel_1_9;
      line_videoOut_rData_frame_line_pixel_1_10 <= line_videoOut_payload_frame_line_pixel_1_10;
      line_videoOut_rData_frame_line_pixel_1_11 <= line_videoOut_payload_frame_line_pixel_1_11;
      line_videoOut_rData_frame_line_pixel_1_12 <= line_videoOut_payload_frame_line_pixel_1_12;
      line_videoOut_rData_frame_line_pixel_1_13 <= line_videoOut_payload_frame_line_pixel_1_13;
      line_videoOut_rData_frame_line_pixel_1_14 <= line_videoOut_payload_frame_line_pixel_1_14;
      line_videoOut_rData_frame_line_pixel_1_15 <= line_videoOut_payload_frame_line_pixel_1_15;
      line_videoOut_rData_frame_line_endOfLine <= line_videoOut_payload_frame_line_endOfLine;
      line_videoOut_rData_frame_endOfFrame <= line_videoOut_payload_frame_endOfFrame;
      line_videoOut_rData_endOfPack <= line_videoOut_payload_endOfPack;
    end
  end


endmodule

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

//VideoFrameHistory replaced by VideoFrameHistory

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//EventM2sPipes replaced by EventM2sPipes

module VideoFrameHistory (
  input      [7:0]    numberOfInputFrames,
  input      [7:0]    numberOfOutputFrames,
  input               videoIn_valid,
  output reg          videoIn_ready,
  input      [15:0]   videoIn_payload_frame_line_pixel_0,
  input      [15:0]   videoIn_payload_frame_line_pixel_1,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [23:0]   videoOut_payload_frame_line_pixel_0,
  output     [23:0]   videoOut_payload_frame_line_pixel_1,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  reg        [47:0]   tmp_ram_port0;
  wire       [13:0]   tmp_inPixelCnt_valueNext;
  wire       [0:0]    tmp_inPixelCnt_valueNext_1;
  wire       [23:0]   tmp_prevData_0_1;
  wire       [23:0]   tmp_prevData_1;
  wire       [23:0]   tmp_postData_0;
  wire       [23:0]   tmp_postData_1;
  wire       [7:0]    tmp_frameCnt_valueNext;
  wire       [0:0]    tmp_frameCnt_valueNext_1;
  wire       [13:0]   tmp_outPixelCnt_valueNext;
  wire       [0:0]    tmp_outPixelCnt_valueNext_1;
  wire       [47:0]   tmp_ram_port;
  wire       [7:0]    tmp_packCnt_valueNext;
  wire       [0:0]    tmp_packCnt_valueNext_1;
  wire       [15:0]   inZero_0;
  wire       [15:0]   inZero_1;
  wire       [23:0]   outZero_0;
  wire       [23:0]   outZero_1;
  wire                videoInPipe_valid;
  wire                videoInPipe_ready;
  wire       [15:0]   videoInPipe_payload_frame_line_pixel_0;
  wire       [15:0]   videoInPipe_payload_frame_line_pixel_1;
  wire                videoInPipe_payload_frame_line_endOfLine;
  wire                videoInPipe_payload_frame_endOfFrame;
  wire                videoInPipe_payload_endOfPack;
  reg                 videoIn_rValid;
  reg        [15:0]   videoIn_rData_frame_line_pixel_0;
  reg        [15:0]   videoIn_rData_frame_line_pixel_1;
  reg                 videoIn_rData_frame_line_endOfLine;
  reg                 videoIn_rData_frame_endOfFrame;
  reg                 videoIn_rData_endOfPack;
  wire                when_Stream_l342;
  reg                 inPixelCnt_willIncrement;
  reg                 inPixelCnt_willClear;
  reg        [13:0]   inPixelCnt_valueNext;
  reg        [13:0]   inPixelCnt_value;
  wire                inPixelCnt_willOverflowIfInc;
  wire                inPixelCnt_willOverflow;
  wire                videoIn_fire;
  wire                when_VideoFrameHistory_l39;
  reg                 firstFrame;
  wire                videoInPipeFire;
  wire                when_VideoFrameHistory_l43;
  wire                when_VideoFrameHistory_l44;
  wire       [47:0]   tmp_prevData_0;
  wire       [23:0]   prevData_0;
  wire       [23:0]   prevData_1;
  wire       [23:0]   postData_0;
  wire       [23:0]   postData_1;
  wire                bridge_valid;
  reg                 bridge_ready;
  wire       [23:0]   bridge_payload_frame_line_pixel_0;
  wire       [23:0]   bridge_payload_frame_line_pixel_1;
  wire                bridge_payload_frame_line_endOfLine;
  wire                bridge_payload_frame_endOfFrame;
  wire                bridge_payload_endOfPack;
  wire                bridgePipe_valid;
  reg                 bridgePipe_ready;
  wire       [23:0]   bridgePipe_payload_frame_line_pixel_0;
  wire       [23:0]   bridgePipe_payload_frame_line_pixel_1;
  wire                bridgePipe_payload_frame_line_endOfLine;
  wire                bridgePipe_payload_frame_endOfFrame;
  wire                bridgePipe_payload_endOfPack;
  reg                 bridge_rValid;
  reg        [23:0]   bridge_rData_frame_line_pixel_0;
  reg        [23:0]   bridge_rData_frame_line_pixel_1;
  reg                 bridge_rData_frame_line_endOfLine;
  reg                 bridge_rData_frame_endOfFrame;
  reg                 bridge_rData_endOfPack;
  wire                when_Stream_l342_1;
  wire                bridgePipeFire;
  reg                 frameCnt_willIncrement;
  reg                 frameCnt_willClear;
  reg        [7:0]    frameCnt_valueNext;
  reg        [7:0]    frameCnt_value;
  wire                frameCnt_willOverflowIfInc;
  wire                frameCnt_willOverflow;
  wire                lastFrame;
  wire                when_VideoFrameHistory_l61;
  wire                when_VideoFrameHistory_l62;
  reg                 outPixelCnt_willIncrement;
  reg                 outPixelCnt_willClear;
  reg        [13:0]   outPixelCnt_valueNext;
  reg        [13:0]   outPixelCnt_value;
  wire                outPixelCnt_willOverflowIfInc;
  wire                outPixelCnt_willOverflow;
  wire                when_VideoFrameHistory_l66;
  reg                 packCnt_willIncrement;
  reg                 packCnt_willClear;
  reg        [7:0]    packCnt_valueNext;
  reg        [7:0]    packCnt_value;
  wire                packCnt_willOverflowIfInc;
  wire                packCnt_willOverflow;
  wire                lastPack;
  wire                when_VideoFrameHistory_l71;
  wire                when_VideoFrameHistory_l72;
  wire                when_Stream_l408;
  reg                 bridgePipe_thrown_valid;
  wire                bridgePipe_thrown_ready;
  wire       [23:0]   bridgePipe_thrown_payload_frame_line_pixel_0;
  wire       [23:0]   bridgePipe_thrown_payload_frame_line_pixel_1;
  wire                bridgePipe_thrown_payload_frame_line_endOfLine;
  wire                bridgePipe_thrown_payload_frame_endOfFrame;
  wire                bridgePipe_thrown_payload_endOfPack;
  reg [47:0] ram [0:16383];

  assign tmp_inPixelCnt_valueNext_1 = inPixelCnt_willIncrement;
  assign tmp_inPixelCnt_valueNext = {13'd0, tmp_inPixelCnt_valueNext_1};
  assign tmp_prevData_0_1 = tmp_prevData_0[23 : 0];
  assign tmp_prevData_1 = tmp_prevData_0[47 : 24];
  assign tmp_postData_0 = {{8{videoInPipe_payload_frame_line_pixel_0[15]}}, videoInPipe_payload_frame_line_pixel_0};
  assign tmp_postData_1 = {{8{videoInPipe_payload_frame_line_pixel_1[15]}}, videoInPipe_payload_frame_line_pixel_1};
  assign tmp_frameCnt_valueNext_1 = frameCnt_willIncrement;
  assign tmp_frameCnt_valueNext = {7'd0, tmp_frameCnt_valueNext_1};
  assign tmp_outPixelCnt_valueNext_1 = outPixelCnt_willIncrement;
  assign tmp_outPixelCnt_valueNext = {13'd0, tmp_outPixelCnt_valueNext_1};
  assign tmp_packCnt_valueNext_1 = packCnt_willIncrement;
  assign tmp_packCnt_valueNext = {7'd0, tmp_packCnt_valueNext_1};
  assign tmp_ram_port = {bridgePipe_payload_frame_line_pixel_1,bridgePipe_payload_frame_line_pixel_0};
  always @(posedge clk) begin
    if(videoIn_ready) begin
      tmp_ram_port0 <= ram[inPixelCnt_value];
    end
  end

  always @(posedge clk) begin
    if(bridgePipeFire) begin
      ram[outPixelCnt_value] <= tmp_ram_port;
    end
  end

  assign inZero_0 = 16'h0;
  assign inZero_1 = 16'h0;
  assign outZero_0 = 24'h0;
  assign outZero_1 = 24'h0;
  always @(*) begin
    videoIn_ready = videoInPipe_ready;
    if(when_Stream_l342) begin
      videoIn_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! videoInPipe_valid);
  assign videoInPipe_valid = videoIn_rValid;
  assign videoInPipe_payload_frame_line_pixel_0 = videoIn_rData_frame_line_pixel_0;
  assign videoInPipe_payload_frame_line_pixel_1 = videoIn_rData_frame_line_pixel_1;
  assign videoInPipe_payload_frame_line_endOfLine = videoIn_rData_frame_line_endOfLine;
  assign videoInPipe_payload_frame_endOfFrame = videoIn_rData_frame_endOfFrame;
  assign videoInPipe_payload_endOfPack = videoIn_rData_endOfPack;
  always @(*) begin
    inPixelCnt_willIncrement = 1'b0;
    if(videoIn_fire) begin
      inPixelCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    inPixelCnt_willClear = 1'b0;
    if(when_VideoFrameHistory_l39) begin
      inPixelCnt_willClear = 1'b1;
    end
  end

  assign inPixelCnt_willOverflowIfInc = (inPixelCnt_value == 14'h3fff);
  assign inPixelCnt_willOverflow = (inPixelCnt_willOverflowIfInc && inPixelCnt_willIncrement);
  always @(*) begin
    inPixelCnt_valueNext = (inPixelCnt_value + tmp_inPixelCnt_valueNext);
    if(inPixelCnt_willClear) begin
      inPixelCnt_valueNext = 14'h0;
    end
  end

  assign videoIn_fire = (videoIn_valid && videoIn_ready);
  assign when_VideoFrameHistory_l39 = (inPixelCnt_willIncrement && videoIn_payload_frame_endOfFrame);
  assign videoInPipeFire = (videoInPipe_valid && videoInPipe_ready);
  assign when_VideoFrameHistory_l43 = (videoInPipe_payload_frame_endOfFrame && videoInPipeFire);
  assign when_VideoFrameHistory_l44 = (videoInPipe_payload_endOfPack && videoInPipeFire);
  assign tmp_prevData_0 = tmp_ram_port0;
  assign prevData_0 = (firstFrame ? outZero_0 : tmp_prevData_0_1);
  assign prevData_1 = (firstFrame ? outZero_1 : tmp_prevData_1);
  assign postData_0 = ($signed(tmp_postData_0) + $signed(prevData_0));
  assign postData_1 = ($signed(tmp_postData_1) + $signed(prevData_1));
  always @(*) begin
    bridge_ready = bridgePipe_ready;
    if(when_Stream_l342_1) begin
      bridge_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! bridgePipe_valid);
  assign bridgePipe_valid = bridge_rValid;
  assign bridgePipe_payload_frame_line_pixel_0 = bridge_rData_frame_line_pixel_0;
  assign bridgePipe_payload_frame_line_pixel_1 = bridge_rData_frame_line_pixel_1;
  assign bridgePipe_payload_frame_line_endOfLine = bridge_rData_frame_line_endOfLine;
  assign bridgePipe_payload_frame_endOfFrame = bridge_rData_frame_endOfFrame;
  assign bridgePipe_payload_endOfPack = bridge_rData_endOfPack;
  assign bridgePipeFire = (bridgePipe_valid && bridgePipe_ready);
  assign bridge_valid = videoInPipe_valid;
  assign videoInPipe_ready = bridge_ready;
  assign bridge_payload_endOfPack = videoInPipe_payload_endOfPack;
  assign bridge_payload_frame_endOfFrame = videoInPipe_payload_frame_endOfFrame;
  assign bridge_payload_frame_line_endOfLine = videoInPipe_payload_frame_line_endOfLine;
  assign bridge_payload_frame_line_pixel_0 = postData_0;
  assign bridge_payload_frame_line_pixel_1 = postData_1;
  always @(*) begin
    frameCnt_willIncrement = 1'b0;
    if(when_VideoFrameHistory_l61) begin
      frameCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    frameCnt_willClear = 1'b0;
    if(when_VideoFrameHistory_l62) begin
      frameCnt_willClear = 1'b1;
    end
  end

  assign frameCnt_willOverflowIfInc = (frameCnt_value == 8'hff);
  assign frameCnt_willOverflow = (frameCnt_willOverflowIfInc && frameCnt_willIncrement);
  always @(*) begin
    frameCnt_valueNext = (frameCnt_value + tmp_frameCnt_valueNext);
    if(frameCnt_willClear) begin
      frameCnt_valueNext = 8'h0;
    end
  end

  assign lastFrame = (frameCnt_value == numberOfInputFrames);
  assign when_VideoFrameHistory_l61 = (bridgePipeFire && bridgePipe_payload_frame_endOfFrame);
  assign when_VideoFrameHistory_l62 = (frameCnt_willIncrement && lastFrame);
  always @(*) begin
    outPixelCnt_willIncrement = 1'b0;
    if(bridgePipeFire) begin
      outPixelCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    outPixelCnt_willClear = 1'b0;
    if(when_VideoFrameHistory_l66) begin
      outPixelCnt_willClear = 1'b1;
    end
  end

  assign outPixelCnt_willOverflowIfInc = (outPixelCnt_value == 14'h3fff);
  assign outPixelCnt_willOverflow = (outPixelCnt_willOverflowIfInc && outPixelCnt_willIncrement);
  always @(*) begin
    outPixelCnt_valueNext = (outPixelCnt_value + tmp_outPixelCnt_valueNext);
    if(outPixelCnt_willClear) begin
      outPixelCnt_valueNext = 14'h0;
    end
  end

  assign when_VideoFrameHistory_l66 = (outPixelCnt_willIncrement && bridgePipe_payload_frame_endOfFrame);
  always @(*) begin
    packCnt_willIncrement = 1'b0;
    if(when_VideoFrameHistory_l71) begin
      packCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    packCnt_willClear = 1'b0;
    if(when_VideoFrameHistory_l72) begin
      packCnt_willClear = 1'b1;
    end
  end

  assign packCnt_willOverflowIfInc = (packCnt_value == 8'hff);
  assign packCnt_willOverflow = (packCnt_willOverflowIfInc && packCnt_willIncrement);
  always @(*) begin
    packCnt_valueNext = (packCnt_value + tmp_packCnt_valueNext);
    if(packCnt_willClear) begin
      packCnt_valueNext = 8'h0;
    end
  end

  assign lastPack = (packCnt_value == numberOfOutputFrames);
  assign when_VideoFrameHistory_l71 = (bridgePipeFire && bridgePipe_payload_endOfPack);
  assign when_VideoFrameHistory_l72 = (packCnt_willIncrement && lastPack);
  assign when_Stream_l408 = (! lastFrame);
  always @(*) begin
    bridgePipe_thrown_valid = bridgePipe_valid;
    if(when_Stream_l408) begin
      bridgePipe_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    bridgePipe_ready = bridgePipe_thrown_ready;
    if(when_Stream_l408) begin
      bridgePipe_ready = 1'b1;
    end
  end

  assign bridgePipe_thrown_payload_frame_line_pixel_0 = bridgePipe_payload_frame_line_pixel_0;
  assign bridgePipe_thrown_payload_frame_line_pixel_1 = bridgePipe_payload_frame_line_pixel_1;
  assign bridgePipe_thrown_payload_frame_line_endOfLine = bridgePipe_payload_frame_line_endOfLine;
  assign bridgePipe_thrown_payload_frame_endOfFrame = bridgePipe_payload_frame_endOfFrame;
  assign bridgePipe_thrown_payload_endOfPack = bridgePipe_payload_endOfPack;
  assign videoOut_valid = bridgePipe_thrown_valid;
  assign bridgePipe_thrown_ready = videoOut_ready;
  assign videoOut_payload_endOfPack = (bridgePipe_payload_endOfPack && lastPack);
  assign videoOut_payload_frame_endOfFrame = bridgePipe_payload_frame_endOfFrame;
  assign videoOut_payload_frame_line_endOfLine = bridgePipe_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_line_pixel_0 = bridgePipe_payload_frame_line_pixel_0;
  assign videoOut_payload_frame_line_pixel_1 = bridgePipe_payload_frame_line_pixel_1;
  always @(posedge clk) begin
    if(reset) begin
      videoIn_rValid <= 1'b0;
      inPixelCnt_value <= 14'h0;
      firstFrame <= 1'b1;
      bridge_rValid <= 1'b0;
      frameCnt_value <= 8'h0;
      outPixelCnt_value <= 14'h0;
      packCnt_value <= 8'h0;
    end else begin
      if(videoIn_ready) begin
        videoIn_rValid <= videoIn_valid;
      end
      inPixelCnt_value <= inPixelCnt_valueNext;
      if(when_VideoFrameHistory_l43) begin
        firstFrame <= 1'b0;
      end
      if(when_VideoFrameHistory_l44) begin
        firstFrame <= 1'b1;
      end
      if(bridge_ready) begin
        bridge_rValid <= bridge_valid;
      end
      frameCnt_value <= frameCnt_valueNext;
      outPixelCnt_value <= outPixelCnt_valueNext;
      packCnt_value <= packCnt_valueNext;
    end
  end

  always @(posedge clk) begin
    if(videoIn_ready) begin
      videoIn_rData_frame_line_pixel_0 <= videoIn_payload_frame_line_pixel_0;
      videoIn_rData_frame_line_pixel_1 <= videoIn_payload_frame_line_pixel_1;
      videoIn_rData_frame_line_endOfLine <= videoIn_payload_frame_line_endOfLine;
      videoIn_rData_frame_endOfFrame <= videoIn_payload_frame_endOfFrame;
      videoIn_rData_endOfPack <= videoIn_payload_endOfPack;
    end
    if(bridge_ready) begin
      bridge_rData_frame_line_pixel_0 <= bridge_payload_frame_line_pixel_0;
      bridge_rData_frame_line_pixel_1 <= bridge_payload_frame_line_pixel_1;
      bridge_rData_frame_line_endOfLine <= bridge_payload_frame_line_endOfLine;
      bridge_rData_frame_endOfFrame <= bridge_payload_frame_endOfFrame;
      bridge_rData_endOfPack <= bridge_payload_endOfPack;
    end
  end


endmodule

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

//SIMD2INT8 replaced by SIMD2INT8

module SIMD2INT8 (
  input      [7:0]    a,
  input      [7:0]    b,
  input      [7:0]    c,
  output     [15:0]   ab,
  output     [15:0]   ac,
  input               CEs_0,
  input               CEs_1,
  input               CEs_2,
  input               CEs_3,
  input               clk
);

  wire       [29:0]   mult_A;
  wire       [17:0]   mult_B;
  wire       [26:0]   mult_D;
  wire       [47:0]   mult_P;
  wire       [29:0]   tmp_A;
  wire       [17:0]   tmp_B;
  wire       [28:0]   tmp_ac_1;
  wire       [15:0]   tmp_ac;
  wire       [15:0]   tmp_ac_2;
  wire       [15:0]   ab_1;
  wire       [15:0]   ac_1;

  assign tmp_A = {{22{b[7]}}, b};
  assign tmp_B = {{10{a[7]}}, a};
  assign tmp_ac_1 = mult_P[47 : 19];
  assign tmp_ac = ($signed(ac_1) + $signed(tmp_ac_2));
  assign tmp_ac_2 = 16'h0001;
  APlusDMultB mult (
    .A        (mult_A[29:0]  ), //i
    .B        (mult_B[17:0]  ), //i
    .D        (mult_D[26:0]  ), //i
    .P        (mult_P[47:0]  ), //o
    .CEs_0    (CEs_0         ), //i
    .CEs_1    (CEs_1         ), //i
    .CEs_2    (CEs_2         ), //i
    .CEs_3    (CEs_3         ), //i
    .clk      (clk           )  //i
  );
  assign mult_A = tmp_A;
  assign mult_D = {c,19'h0};
  assign mult_B = tmp_B;
  assign ab_1 = mult_P[15 : 0];
  assign ac_1 = tmp_ac_1[15 : 0];
  assign ab = ab_1;
  assign ac = (ab_1[15] ? tmp_ac : ac_1);

endmodule

module EventM2sPipes (
  input               eventIn_valid,
  output              eventIn_ready,
  output              eventOut_valid,
  input               eventOut_ready,
  output              CEs_0,
  output              CEs_1,
  output              CEs_2,
  output              CEs_3,
  output              CEs_4,
  output              CEs_5,
  output              CEs_6,
  output              CEs_7,
  output              CEs_8,
  input               clk,
  input               reset
);

  wire                events_0_valid;
  reg                 events_0_ready;
  wire                events_1_valid;
  reg                 events_1_ready;
  wire                events_2_valid;
  reg                 events_2_ready;
  wire                events_3_valid;
  reg                 events_3_ready;
  wire                events_4_valid;
  reg                 events_4_ready;
  wire                events_5_valid;
  reg                 events_5_ready;
  wire                events_6_valid;
  reg                 events_6_ready;
  wire                events_7_valid;
  reg                 events_7_ready;
  wire                events_8_valid;
  reg                 events_8_ready;
  wire                events_0_m2sPipe_valid;
  wire                events_0_m2sPipe_ready;
  reg                 events_0_rValid;
  wire                when_Stream_l342;
  wire                events_1_m2sPipe_valid;
  wire                events_1_m2sPipe_ready;
  reg                 events_1_rValid;
  wire                when_Stream_l342_1;
  wire                events_2_m2sPipe_valid;
  wire                events_2_m2sPipe_ready;
  reg                 events_2_rValid;
  wire                when_Stream_l342_2;
  wire                events_3_m2sPipe_valid;
  wire                events_3_m2sPipe_ready;
  reg                 events_3_rValid;
  wire                when_Stream_l342_3;
  wire                events_4_m2sPipe_valid;
  wire                events_4_m2sPipe_ready;
  reg                 events_4_rValid;
  wire                when_Stream_l342_4;
  wire                events_5_m2sPipe_valid;
  wire                events_5_m2sPipe_ready;
  reg                 events_5_rValid;
  wire                when_Stream_l342_5;
  wire                events_6_m2sPipe_valid;
  wire                events_6_m2sPipe_ready;
  reg                 events_6_rValid;
  wire                when_Stream_l342_6;
  wire                events_7_m2sPipe_valid;
  wire                events_7_m2sPipe_ready;
  reg                 events_7_rValid;
  wire                when_Stream_l342_7;
  wire                events_8_m2sPipe_valid;
  wire                events_8_m2sPipe_ready;
  reg                 events_8_rValid;
  wire                when_Stream_l342_8;

  assign CEs_0 = events_0_ready;
  assign CEs_1 = events_1_ready;
  assign CEs_2 = events_2_ready;
  assign CEs_3 = events_3_ready;
  assign CEs_4 = events_4_ready;
  assign CEs_5 = events_5_ready;
  assign CEs_6 = events_6_ready;
  assign CEs_7 = events_7_ready;
  assign CEs_8 = events_8_ready;
  assign events_0_valid = eventIn_valid;
  assign eventIn_ready = events_0_ready;
  always @(*) begin
    events_0_ready = events_0_m2sPipe_ready;
    if(when_Stream_l342) begin
      events_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! events_0_m2sPipe_valid);
  assign events_0_m2sPipe_valid = events_0_rValid;
  assign events_1_valid = events_0_m2sPipe_valid;
  assign events_0_m2sPipe_ready = events_1_ready;
  always @(*) begin
    events_1_ready = events_1_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      events_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! events_1_m2sPipe_valid);
  assign events_1_m2sPipe_valid = events_1_rValid;
  assign events_2_valid = events_1_m2sPipe_valid;
  assign events_1_m2sPipe_ready = events_2_ready;
  always @(*) begin
    events_2_ready = events_2_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      events_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! events_2_m2sPipe_valid);
  assign events_2_m2sPipe_valid = events_2_rValid;
  assign events_3_valid = events_2_m2sPipe_valid;
  assign events_2_m2sPipe_ready = events_3_ready;
  always @(*) begin
    events_3_ready = events_3_m2sPipe_ready;
    if(when_Stream_l342_3) begin
      events_3_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! events_3_m2sPipe_valid);
  assign events_3_m2sPipe_valid = events_3_rValid;
  assign events_4_valid = events_3_m2sPipe_valid;
  assign events_3_m2sPipe_ready = events_4_ready;
  always @(*) begin
    events_4_ready = events_4_m2sPipe_ready;
    if(when_Stream_l342_4) begin
      events_4_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! events_4_m2sPipe_valid);
  assign events_4_m2sPipe_valid = events_4_rValid;
  assign events_5_valid = events_4_m2sPipe_valid;
  assign events_4_m2sPipe_ready = events_5_ready;
  always @(*) begin
    events_5_ready = events_5_m2sPipe_ready;
    if(when_Stream_l342_5) begin
      events_5_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! events_5_m2sPipe_valid);
  assign events_5_m2sPipe_valid = events_5_rValid;
  assign events_6_valid = events_5_m2sPipe_valid;
  assign events_5_m2sPipe_ready = events_6_ready;
  always @(*) begin
    events_6_ready = events_6_m2sPipe_ready;
    if(when_Stream_l342_6) begin
      events_6_ready = 1'b1;
    end
  end

  assign when_Stream_l342_6 = (! events_6_m2sPipe_valid);
  assign events_6_m2sPipe_valid = events_6_rValid;
  assign events_7_valid = events_6_m2sPipe_valid;
  assign events_6_m2sPipe_ready = events_7_ready;
  always @(*) begin
    events_7_ready = events_7_m2sPipe_ready;
    if(when_Stream_l342_7) begin
      events_7_ready = 1'b1;
    end
  end

  assign when_Stream_l342_7 = (! events_7_m2sPipe_valid);
  assign events_7_m2sPipe_valid = events_7_rValid;
  assign events_8_valid = events_7_m2sPipe_valid;
  assign events_7_m2sPipe_ready = events_8_ready;
  always @(*) begin
    events_8_ready = events_8_m2sPipe_ready;
    if(when_Stream_l342_8) begin
      events_8_ready = 1'b1;
    end
  end

  assign when_Stream_l342_8 = (! events_8_m2sPipe_valid);
  assign events_8_m2sPipe_valid = events_8_rValid;
  assign eventOut_valid = events_8_m2sPipe_valid;
  assign events_8_m2sPipe_ready = eventOut_ready;
  always @(posedge clk) begin
    if(reset) begin
      events_0_rValid <= 1'b0;
      events_1_rValid <= 1'b0;
      events_2_rValid <= 1'b0;
      events_3_rValid <= 1'b0;
      events_4_rValid <= 1'b0;
      events_5_rValid <= 1'b0;
      events_6_rValid <= 1'b0;
      events_7_rValid <= 1'b0;
      events_8_rValid <= 1'b0;
    end else begin
      if(events_0_ready) begin
        events_0_rValid <= events_0_valid;
      end
      if(events_1_ready) begin
        events_1_rValid <= events_1_valid;
      end
      if(events_2_ready) begin
        events_2_rValid <= events_2_valid;
      end
      if(events_3_ready) begin
        events_3_rValid <= events_3_valid;
      end
      if(events_4_ready) begin
        events_4_rValid <= events_4_valid;
      end
      if(events_5_ready) begin
        events_5_rValid <= events_5_valid;
      end
      if(events_6_ready) begin
        events_6_rValid <= events_6_valid;
      end
      if(events_7_ready) begin
        events_7_rValid <= events_7_valid;
      end
      if(events_8_ready) begin
        events_8_rValid <= events_8_valid;
      end
    end
  end


endmodule

module PixelBufferSame (
  input               videoIn_valid,
  output reg          videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_15,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_15,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_2_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  wire       [7:0]    tmp_pixelBuffer;
  wire       [87:0]   tmp_pixelBuffer_1;
  wire       [7:0]    tmp_pixelBuffer_2;
  wire       [39:0]   tmp_pixelBuffer_3;
  wire       [7:0]    tmp_pixelBuffer_4;
  wire       [95:0]   tmp_pixelBuffer_5;
  wire       [7:0]    tmp_pixelBuffer_6;
  wire       [47:0]   tmp_pixelBuffer_7;
  wire       [7:0]    tmp_pixelBuffer_8;
  wire       [95:0]   tmp_pixelBuffer_9;
  wire       [7:0]    tmp_pixelBuffer_10;
  wire       [47:0]   tmp_pixelBuffer_11;
  wire       [383:0]  tmp_pixelBuffer_12;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0;
  wire       [87:0]   tmp_tmp_pixelVec_0_0_0_1;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_2;
  wire       [39:0]   tmp_tmp_pixelVec_0_0_0_3;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_4;
  wire       [95:0]   tmp_tmp_pixelVec_0_0_0_5;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_6;
  wire       [47:0]   tmp_tmp_pixelVec_0_0_0_7;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_8;
  wire       [95:0]   tmp_tmp_pixelVec_0_0_0_9;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_10;
  wire       [47:0]   tmp_tmp_pixelVec_0_0_0_11;
  wire       [7:0]    zero_0_0;
  wire       [7:0]    zero_0_1;
  wire       [7:0]    zero_0_2;
  wire       [7:0]    zero_0_3;
  wire       [7:0]    zero_0_4;
  wire       [7:0]    zero_0_5;
  wire       [7:0]    zero_0_6;
  wire       [7:0]    zero_0_7;
  wire       [7:0]    zero_0_8;
  wire       [7:0]    zero_0_9;
  wire       [7:0]    zero_0_10;
  wire       [7:0]    zero_0_11;
  wire       [7:0]    zero_0_12;
  wire       [7:0]    zero_0_13;
  wire       [7:0]    zero_0_14;
  wire       [7:0]    zero_0_15;
  wire       [7:0]    zero_1_0;
  wire       [7:0]    zero_1_1;
  wire       [7:0]    zero_1_2;
  wire       [7:0]    zero_1_3;
  wire       [7:0]    zero_1_4;
  wire       [7:0]    zero_1_5;
  wire       [7:0]    zero_1_6;
  wire       [7:0]    zero_1_7;
  wire       [7:0]    zero_1_8;
  wire       [7:0]    zero_1_9;
  wire       [7:0]    zero_1_10;
  wire       [7:0]    zero_1_11;
  wire       [7:0]    zero_1_12;
  wire       [7:0]    zero_1_13;
  wire       [7:0]    zero_1_14;
  wire       [7:0]    zero_1_15;
  wire       [7:0]    zero_2_0;
  wire       [7:0]    zero_2_1;
  wire       [7:0]    zero_2_2;
  wire       [7:0]    zero_2_3;
  wire       [7:0]    zero_2_4;
  wire       [7:0]    zero_2_5;
  wire       [7:0]    zero_2_6;
  wire       [7:0]    zero_2_7;
  wire       [7:0]    zero_2_8;
  wire       [7:0]    zero_2_9;
  wire       [7:0]    zero_2_10;
  wire       [7:0]    zero_2_11;
  wire       [7:0]    zero_2_12;
  wire       [7:0]    zero_2_13;
  wire       [7:0]    zero_2_14;
  wire       [7:0]    zero_2_15;
  wire       [383:0]  tmp_zero_0_0;
  wire       [127:0]  tmp_zero_0_0_1;
  wire       [127:0]  tmp_zero_1_0;
  wire       [127:0]  tmp_zero_2_0;
  wire                padded_valid;
  wire                padded_ready;
  wire       [7:0]    padded_payload_frame_line_pixel_0_0;
  wire       [7:0]    padded_payload_frame_line_pixel_0_1;
  wire       [7:0]    padded_payload_frame_line_pixel_0_2;
  wire       [7:0]    padded_payload_frame_line_pixel_0_3;
  wire       [7:0]    padded_payload_frame_line_pixel_0_4;
  wire       [7:0]    padded_payload_frame_line_pixel_0_5;
  wire       [7:0]    padded_payload_frame_line_pixel_0_6;
  wire       [7:0]    padded_payload_frame_line_pixel_0_7;
  wire       [7:0]    padded_payload_frame_line_pixel_0_8;
  wire       [7:0]    padded_payload_frame_line_pixel_0_9;
  wire       [7:0]    padded_payload_frame_line_pixel_0_10;
  wire       [7:0]    padded_payload_frame_line_pixel_0_11;
  wire       [7:0]    padded_payload_frame_line_pixel_0_12;
  wire       [7:0]    padded_payload_frame_line_pixel_0_13;
  wire       [7:0]    padded_payload_frame_line_pixel_0_14;
  wire       [7:0]    padded_payload_frame_line_pixel_0_15;
  wire       [7:0]    padded_payload_frame_line_pixel_1_0;
  wire       [7:0]    padded_payload_frame_line_pixel_1_1;
  wire       [7:0]    padded_payload_frame_line_pixel_1_2;
  wire       [7:0]    padded_payload_frame_line_pixel_1_3;
  wire       [7:0]    padded_payload_frame_line_pixel_1_4;
  wire       [7:0]    padded_payload_frame_line_pixel_1_5;
  wire       [7:0]    padded_payload_frame_line_pixel_1_6;
  wire       [7:0]    padded_payload_frame_line_pixel_1_7;
  wire       [7:0]    padded_payload_frame_line_pixel_1_8;
  wire       [7:0]    padded_payload_frame_line_pixel_1_9;
  wire       [7:0]    padded_payload_frame_line_pixel_1_10;
  wire       [7:0]    padded_payload_frame_line_pixel_1_11;
  wire       [7:0]    padded_payload_frame_line_pixel_1_12;
  wire       [7:0]    padded_payload_frame_line_pixel_1_13;
  wire       [7:0]    padded_payload_frame_line_pixel_1_14;
  wire       [7:0]    padded_payload_frame_line_pixel_1_15;
  wire       [7:0]    padded_payload_frame_line_pixel_2_0;
  wire       [7:0]    padded_payload_frame_line_pixel_2_1;
  wire       [7:0]    padded_payload_frame_line_pixel_2_2;
  wire       [7:0]    padded_payload_frame_line_pixel_2_3;
  wire       [7:0]    padded_payload_frame_line_pixel_2_4;
  wire       [7:0]    padded_payload_frame_line_pixel_2_5;
  wire       [7:0]    padded_payload_frame_line_pixel_2_6;
  wire       [7:0]    padded_payload_frame_line_pixel_2_7;
  wire       [7:0]    padded_payload_frame_line_pixel_2_8;
  wire       [7:0]    padded_payload_frame_line_pixel_2_9;
  wire       [7:0]    padded_payload_frame_line_pixel_2_10;
  wire       [7:0]    padded_payload_frame_line_pixel_2_11;
  wire       [7:0]    padded_payload_frame_line_pixel_2_12;
  wire       [7:0]    padded_payload_frame_line_pixel_2_13;
  wire       [7:0]    padded_payload_frame_line_pixel_2_14;
  wire       [7:0]    padded_payload_frame_line_pixel_2_15;
  wire                padded_payload_frame_line_endOfLine;
  wire                padded_payload_frame_endOfFrame;
  wire                padded_payload_endOfPack;
  wire                videoInFire;
  wire                videoOutFire;
  wire                paddedFire;
  wire                when_PixelBufferSame_l46;
  reg                 tmp_bridge_payload_endOfPack;
  wire                tmp_bridge_payload_endOfPack_1;
  wire                tmp_bridge_payload_endOfPack_2;
  reg                 paddedCond;
  wire                when_PixelBufferSame_l48;
  reg                 tmp_padded_valid;
  reg        [767:0]  pixelBuffer;
  wire                bridge_valid;
  reg                 bridge_ready;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_2_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_2_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_0_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_1_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_2_2_15;
  wire                bridge_payload_frame_line_endOfLine;
  wire                bridge_payload_frame_endOfFrame;
  wire                bridge_payload_endOfPack;
  wire                bridgeFire;
  reg        [1:0]    cntPrev;
  reg        [1:0]    cntPost;
  wire                cntPrevStable;
  wire                cntPostStable;
  wire                cntPrevEqualVec_0;
  wire                cntPostEqualVec_0;
  wire                when_PixelBufferSame_l74;
  wire                when_PixelBufferSame_l75;
  wire                when_PixelBufferSame_l76;
  wire                when_PixelBufferSame_l77;
  wire       [7:0]    pixelVec_0_0_0;
  wire       [7:0]    pixelVec_0_0_1;
  wire       [7:0]    pixelVec_0_0_2;
  wire       [7:0]    pixelVec_0_0_3;
  wire       [7:0]    pixelVec_0_0_4;
  wire       [7:0]    pixelVec_0_0_5;
  wire       [7:0]    pixelVec_0_0_6;
  wire       [7:0]    pixelVec_0_0_7;
  wire       [7:0]    pixelVec_0_0_8;
  wire       [7:0]    pixelVec_0_0_9;
  wire       [7:0]    pixelVec_0_0_10;
  wire       [7:0]    pixelVec_0_0_11;
  wire       [7:0]    pixelVec_0_0_12;
  wire       [7:0]    pixelVec_0_0_13;
  wire       [7:0]    pixelVec_0_0_14;
  wire       [7:0]    pixelVec_0_0_15;
  wire       [7:0]    pixelVec_0_1_0;
  wire       [7:0]    pixelVec_0_1_1;
  wire       [7:0]    pixelVec_0_1_2;
  wire       [7:0]    pixelVec_0_1_3;
  wire       [7:0]    pixelVec_0_1_4;
  wire       [7:0]    pixelVec_0_1_5;
  wire       [7:0]    pixelVec_0_1_6;
  wire       [7:0]    pixelVec_0_1_7;
  wire       [7:0]    pixelVec_0_1_8;
  wire       [7:0]    pixelVec_0_1_9;
  wire       [7:0]    pixelVec_0_1_10;
  wire       [7:0]    pixelVec_0_1_11;
  wire       [7:0]    pixelVec_0_1_12;
  wire       [7:0]    pixelVec_0_1_13;
  wire       [7:0]    pixelVec_0_1_14;
  wire       [7:0]    pixelVec_0_1_15;
  wire       [7:0]    pixelVec_0_2_0;
  wire       [7:0]    pixelVec_0_2_1;
  wire       [7:0]    pixelVec_0_2_2;
  wire       [7:0]    pixelVec_0_2_3;
  wire       [7:0]    pixelVec_0_2_4;
  wire       [7:0]    pixelVec_0_2_5;
  wire       [7:0]    pixelVec_0_2_6;
  wire       [7:0]    pixelVec_0_2_7;
  wire       [7:0]    pixelVec_0_2_8;
  wire       [7:0]    pixelVec_0_2_9;
  wire       [7:0]    pixelVec_0_2_10;
  wire       [7:0]    pixelVec_0_2_11;
  wire       [7:0]    pixelVec_0_2_12;
  wire       [7:0]    pixelVec_0_2_13;
  wire       [7:0]    pixelVec_0_2_14;
  wire       [7:0]    pixelVec_0_2_15;
  wire       [7:0]    pixelVec_1_0_0;
  wire       [7:0]    pixelVec_1_0_1;
  wire       [7:0]    pixelVec_1_0_2;
  wire       [7:0]    pixelVec_1_0_3;
  wire       [7:0]    pixelVec_1_0_4;
  wire       [7:0]    pixelVec_1_0_5;
  wire       [7:0]    pixelVec_1_0_6;
  wire       [7:0]    pixelVec_1_0_7;
  wire       [7:0]    pixelVec_1_0_8;
  wire       [7:0]    pixelVec_1_0_9;
  wire       [7:0]    pixelVec_1_0_10;
  wire       [7:0]    pixelVec_1_0_11;
  wire       [7:0]    pixelVec_1_0_12;
  wire       [7:0]    pixelVec_1_0_13;
  wire       [7:0]    pixelVec_1_0_14;
  wire       [7:0]    pixelVec_1_0_15;
  wire       [7:0]    pixelVec_1_1_0;
  wire       [7:0]    pixelVec_1_1_1;
  wire       [7:0]    pixelVec_1_1_2;
  wire       [7:0]    pixelVec_1_1_3;
  wire       [7:0]    pixelVec_1_1_4;
  wire       [7:0]    pixelVec_1_1_5;
  wire       [7:0]    pixelVec_1_1_6;
  wire       [7:0]    pixelVec_1_1_7;
  wire       [7:0]    pixelVec_1_1_8;
  wire       [7:0]    pixelVec_1_1_9;
  wire       [7:0]    pixelVec_1_1_10;
  wire       [7:0]    pixelVec_1_1_11;
  wire       [7:0]    pixelVec_1_1_12;
  wire       [7:0]    pixelVec_1_1_13;
  wire       [7:0]    pixelVec_1_1_14;
  wire       [7:0]    pixelVec_1_1_15;
  wire       [7:0]    pixelVec_1_2_0;
  wire       [7:0]    pixelVec_1_2_1;
  wire       [7:0]    pixelVec_1_2_2;
  wire       [7:0]    pixelVec_1_2_3;
  wire       [7:0]    pixelVec_1_2_4;
  wire       [7:0]    pixelVec_1_2_5;
  wire       [7:0]    pixelVec_1_2_6;
  wire       [7:0]    pixelVec_1_2_7;
  wire       [7:0]    pixelVec_1_2_8;
  wire       [7:0]    pixelVec_1_2_9;
  wire       [7:0]    pixelVec_1_2_10;
  wire       [7:0]    pixelVec_1_2_11;
  wire       [7:0]    pixelVec_1_2_12;
  wire       [7:0]    pixelVec_1_2_13;
  wire       [7:0]    pixelVec_1_2_14;
  wire       [7:0]    pixelVec_1_2_15;
  wire       [7:0]    pixelVec_2_0_0;
  wire       [7:0]    pixelVec_2_0_1;
  wire       [7:0]    pixelVec_2_0_2;
  wire       [7:0]    pixelVec_2_0_3;
  wire       [7:0]    pixelVec_2_0_4;
  wire       [7:0]    pixelVec_2_0_5;
  wire       [7:0]    pixelVec_2_0_6;
  wire       [7:0]    pixelVec_2_0_7;
  wire       [7:0]    pixelVec_2_0_8;
  wire       [7:0]    pixelVec_2_0_9;
  wire       [7:0]    pixelVec_2_0_10;
  wire       [7:0]    pixelVec_2_0_11;
  wire       [7:0]    pixelVec_2_0_12;
  wire       [7:0]    pixelVec_2_0_13;
  wire       [7:0]    pixelVec_2_0_14;
  wire       [7:0]    pixelVec_2_0_15;
  wire       [7:0]    pixelVec_2_1_0;
  wire       [7:0]    pixelVec_2_1_1;
  wire       [7:0]    pixelVec_2_1_2;
  wire       [7:0]    pixelVec_2_1_3;
  wire       [7:0]    pixelVec_2_1_4;
  wire       [7:0]    pixelVec_2_1_5;
  wire       [7:0]    pixelVec_2_1_6;
  wire       [7:0]    pixelVec_2_1_7;
  wire       [7:0]    pixelVec_2_1_8;
  wire       [7:0]    pixelVec_2_1_9;
  wire       [7:0]    pixelVec_2_1_10;
  wire       [7:0]    pixelVec_2_1_11;
  wire       [7:0]    pixelVec_2_1_12;
  wire       [7:0]    pixelVec_2_1_13;
  wire       [7:0]    pixelVec_2_1_14;
  wire       [7:0]    pixelVec_2_1_15;
  wire       [7:0]    pixelVec_2_2_0;
  wire       [7:0]    pixelVec_2_2_1;
  wire       [7:0]    pixelVec_2_2_2;
  wire       [7:0]    pixelVec_2_2_3;
  wire       [7:0]    pixelVec_2_2_4;
  wire       [7:0]    pixelVec_2_2_5;
  wire       [7:0]    pixelVec_2_2_6;
  wire       [7:0]    pixelVec_2_2_7;
  wire       [7:0]    pixelVec_2_2_8;
  wire       [7:0]    pixelVec_2_2_9;
  wire       [7:0]    pixelVec_2_2_10;
  wire       [7:0]    pixelVec_2_2_11;
  wire       [7:0]    pixelVec_2_2_12;
  wire       [7:0]    pixelVec_2_2_13;
  wire       [7:0]    pixelVec_2_2_14;
  wire       [7:0]    pixelVec_2_2_15;
  wire       [1151:0] tmp_pixelVec_0_0_0;
  wire       [383:0]  tmp_pixelVec_0_0_0_1;
  wire       [127:0]  tmp_pixelVec_0_0_0_2;
  wire       [127:0]  tmp_pixelVec_0_1_0;
  wire       [127:0]  tmp_pixelVec_0_2_0;
  wire       [383:0]  tmp_pixelVec_1_0_0;
  wire       [127:0]  tmp_pixelVec_1_0_0_1;
  wire       [127:0]  tmp_pixelVec_1_1_0;
  wire       [127:0]  tmp_pixelVec_1_2_0;
  wire       [383:0]  tmp_pixelVec_2_0_0;
  wire       [127:0]  tmp_pixelVec_2_0_0_1;
  wire       [127:0]  tmp_pixelVec_2_1_0;
  wire       [127:0]  tmp_pixelVec_2_2_0;
  wire       [7:0]    up_0_0_0;
  wire       [7:0]    up_0_0_1;
  wire       [7:0]    up_0_0_2;
  wire       [7:0]    up_0_0_3;
  wire       [7:0]    up_0_0_4;
  wire       [7:0]    up_0_0_5;
  wire       [7:0]    up_0_0_6;
  wire       [7:0]    up_0_0_7;
  wire       [7:0]    up_0_0_8;
  wire       [7:0]    up_0_0_9;
  wire       [7:0]    up_0_0_10;
  wire       [7:0]    up_0_0_11;
  wire       [7:0]    up_0_0_12;
  wire       [7:0]    up_0_0_13;
  wire       [7:0]    up_0_0_14;
  wire       [7:0]    up_0_0_15;
  wire       [7:0]    up_0_1_0;
  wire       [7:0]    up_0_1_1;
  wire       [7:0]    up_0_1_2;
  wire       [7:0]    up_0_1_3;
  wire       [7:0]    up_0_1_4;
  wire       [7:0]    up_0_1_5;
  wire       [7:0]    up_0_1_6;
  wire       [7:0]    up_0_1_7;
  wire       [7:0]    up_0_1_8;
  wire       [7:0]    up_0_1_9;
  wire       [7:0]    up_0_1_10;
  wire       [7:0]    up_0_1_11;
  wire       [7:0]    up_0_1_12;
  wire       [7:0]    up_0_1_13;
  wire       [7:0]    up_0_1_14;
  wire       [7:0]    up_0_1_15;
  wire       [7:0]    up_0_2_0;
  wire       [7:0]    up_0_2_1;
  wire       [7:0]    up_0_2_2;
  wire       [7:0]    up_0_2_3;
  wire       [7:0]    up_0_2_4;
  wire       [7:0]    up_0_2_5;
  wire       [7:0]    up_0_2_6;
  wire       [7:0]    up_0_2_7;
  wire       [7:0]    up_0_2_8;
  wire       [7:0]    up_0_2_9;
  wire       [7:0]    up_0_2_10;
  wire       [7:0]    up_0_2_11;
  wire       [7:0]    up_0_2_12;
  wire       [7:0]    up_0_2_13;
  wire       [7:0]    up_0_2_14;
  wire       [7:0]    up_0_2_15;
  wire       [7:0]    down_0_0_0;
  wire       [7:0]    down_0_0_1;
  wire       [7:0]    down_0_0_2;
  wire       [7:0]    down_0_0_3;
  wire       [7:0]    down_0_0_4;
  wire       [7:0]    down_0_0_5;
  wire       [7:0]    down_0_0_6;
  wire       [7:0]    down_0_0_7;
  wire       [7:0]    down_0_0_8;
  wire       [7:0]    down_0_0_9;
  wire       [7:0]    down_0_0_10;
  wire       [7:0]    down_0_0_11;
  wire       [7:0]    down_0_0_12;
  wire       [7:0]    down_0_0_13;
  wire       [7:0]    down_0_0_14;
  wire       [7:0]    down_0_0_15;
  wire       [7:0]    down_0_1_0;
  wire       [7:0]    down_0_1_1;
  wire       [7:0]    down_0_1_2;
  wire       [7:0]    down_0_1_3;
  wire       [7:0]    down_0_1_4;
  wire       [7:0]    down_0_1_5;
  wire       [7:0]    down_0_1_6;
  wire       [7:0]    down_0_1_7;
  wire       [7:0]    down_0_1_8;
  wire       [7:0]    down_0_1_9;
  wire       [7:0]    down_0_1_10;
  wire       [7:0]    down_0_1_11;
  wire       [7:0]    down_0_1_12;
  wire       [7:0]    down_0_1_13;
  wire       [7:0]    down_0_1_14;
  wire       [7:0]    down_0_1_15;
  wire       [7:0]    down_0_2_0;
  wire       [7:0]    down_0_2_1;
  wire       [7:0]    down_0_2_2;
  wire       [7:0]    down_0_2_3;
  wire       [7:0]    down_0_2_4;
  wire       [7:0]    down_0_2_5;
  wire       [7:0]    down_0_2_6;
  wire       [7:0]    down_0_2_7;
  wire       [7:0]    down_0_2_8;
  wire       [7:0]    down_0_2_9;
  wire       [7:0]    down_0_2_10;
  wire       [7:0]    down_0_2_11;
  wire       [7:0]    down_0_2_12;
  wire       [7:0]    down_0_2_13;
  wire       [7:0]    down_0_2_14;
  wire       [7:0]    down_0_2_15;
  reg                 padded_payload_frame_endOfFrame_delay_1;
  reg                 padded_payload_frame_line_endOfLine_delay_1;
  reg                 cnt_willIncrement;
  reg                 cnt_willClear;
  reg        [0:0]    cnt_valueNext;
  reg        [0:0]    cnt_value;
  wire                cnt_willOverflowIfInc;
  wire                cnt_willOverflow;
  wire                cntWontOverflowIfInc;
  wire                when_PixelBufferSame_l92;
  wire                when_PixelBufferSame_l93;
  reg                 tmp_videoOut_valid;

  assign tmp_pixelBuffer_12 = (pixelBuffer >>> 384);
  assign tmp_pixelBuffer = padded_payload_frame_line_pixel_2_11;
  assign tmp_pixelBuffer_1 = {padded_payload_frame_line_pixel_2_10,{padded_payload_frame_line_pixel_2_9,{padded_payload_frame_line_pixel_2_8,{padded_payload_frame_line_pixel_2_7,{padded_payload_frame_line_pixel_2_6,{tmp_pixelBuffer_2,tmp_pixelBuffer_3}}}}}};
  assign tmp_pixelBuffer_4 = padded_payload_frame_line_pixel_1_12;
  assign tmp_pixelBuffer_5 = {padded_payload_frame_line_pixel_1_11,{padded_payload_frame_line_pixel_1_10,{padded_payload_frame_line_pixel_1_9,{padded_payload_frame_line_pixel_1_8,{padded_payload_frame_line_pixel_1_7,{tmp_pixelBuffer_6,tmp_pixelBuffer_7}}}}}};
  assign tmp_pixelBuffer_8 = padded_payload_frame_line_pixel_0_12;
  assign tmp_pixelBuffer_9 = {padded_payload_frame_line_pixel_0_11,{padded_payload_frame_line_pixel_0_10,{padded_payload_frame_line_pixel_0_9,{padded_payload_frame_line_pixel_0_8,{padded_payload_frame_line_pixel_0_7,{tmp_pixelBuffer_10,tmp_pixelBuffer_11}}}}}};
  assign tmp_pixelBuffer_2 = padded_payload_frame_line_pixel_2_5;
  assign tmp_pixelBuffer_3 = {padded_payload_frame_line_pixel_2_4,{padded_payload_frame_line_pixel_2_3,{padded_payload_frame_line_pixel_2_2,{padded_payload_frame_line_pixel_2_1,padded_payload_frame_line_pixel_2_0}}}};
  assign tmp_pixelBuffer_6 = padded_payload_frame_line_pixel_1_6;
  assign tmp_pixelBuffer_7 = {padded_payload_frame_line_pixel_1_5,{padded_payload_frame_line_pixel_1_4,{padded_payload_frame_line_pixel_1_3,{padded_payload_frame_line_pixel_1_2,{padded_payload_frame_line_pixel_1_1,padded_payload_frame_line_pixel_1_0}}}}};
  assign tmp_pixelBuffer_10 = padded_payload_frame_line_pixel_0_6;
  assign tmp_pixelBuffer_11 = {padded_payload_frame_line_pixel_0_5,{padded_payload_frame_line_pixel_0_4,{padded_payload_frame_line_pixel_0_3,{padded_payload_frame_line_pixel_0_2,{padded_payload_frame_line_pixel_0_1,padded_payload_frame_line_pixel_0_0}}}}};
  assign tmp_tmp_pixelVec_0_0_0 = videoIn_payload_frame_line_pixel_2_11;
  assign tmp_tmp_pixelVec_0_0_0_1 = {videoIn_payload_frame_line_pixel_2_10,{videoIn_payload_frame_line_pixel_2_9,{videoIn_payload_frame_line_pixel_2_8,{videoIn_payload_frame_line_pixel_2_7,{videoIn_payload_frame_line_pixel_2_6,{tmp_tmp_pixelVec_0_0_0_2,tmp_tmp_pixelVec_0_0_0_3}}}}}};
  assign tmp_tmp_pixelVec_0_0_0_4 = videoIn_payload_frame_line_pixel_1_12;
  assign tmp_tmp_pixelVec_0_0_0_5 = {videoIn_payload_frame_line_pixel_1_11,{videoIn_payload_frame_line_pixel_1_10,{videoIn_payload_frame_line_pixel_1_9,{videoIn_payload_frame_line_pixel_1_8,{videoIn_payload_frame_line_pixel_1_7,{tmp_tmp_pixelVec_0_0_0_6,tmp_tmp_pixelVec_0_0_0_7}}}}}};
  assign tmp_tmp_pixelVec_0_0_0_8 = videoIn_payload_frame_line_pixel_0_12;
  assign tmp_tmp_pixelVec_0_0_0_9 = {videoIn_payload_frame_line_pixel_0_11,{videoIn_payload_frame_line_pixel_0_10,{videoIn_payload_frame_line_pixel_0_9,{videoIn_payload_frame_line_pixel_0_8,{videoIn_payload_frame_line_pixel_0_7,{tmp_tmp_pixelVec_0_0_0_10,tmp_tmp_pixelVec_0_0_0_11}}}}}};
  assign tmp_tmp_pixelVec_0_0_0_2 = videoIn_payload_frame_line_pixel_2_5;
  assign tmp_tmp_pixelVec_0_0_0_3 = {videoIn_payload_frame_line_pixel_2_4,{videoIn_payload_frame_line_pixel_2_3,{videoIn_payload_frame_line_pixel_2_2,{videoIn_payload_frame_line_pixel_2_1,videoIn_payload_frame_line_pixel_2_0}}}};
  assign tmp_tmp_pixelVec_0_0_0_6 = videoIn_payload_frame_line_pixel_1_6;
  assign tmp_tmp_pixelVec_0_0_0_7 = {videoIn_payload_frame_line_pixel_1_5,{videoIn_payload_frame_line_pixel_1_4,{videoIn_payload_frame_line_pixel_1_3,{videoIn_payload_frame_line_pixel_1_2,{videoIn_payload_frame_line_pixel_1_1,videoIn_payload_frame_line_pixel_1_0}}}}};
  assign tmp_tmp_pixelVec_0_0_0_10 = videoIn_payload_frame_line_pixel_0_6;
  assign tmp_tmp_pixelVec_0_0_0_11 = {videoIn_payload_frame_line_pixel_0_5,{videoIn_payload_frame_line_pixel_0_4,{videoIn_payload_frame_line_pixel_0_3,{videoIn_payload_frame_line_pixel_0_2,{videoIn_payload_frame_line_pixel_0_1,videoIn_payload_frame_line_pixel_0_0}}}}};
  assign tmp_zero_0_0 = 384'h0;
  assign tmp_zero_0_0_1 = tmp_zero_0_0[127 : 0];
  assign zero_0_0 = tmp_zero_0_0_1[7 : 0];
  assign zero_0_1 = tmp_zero_0_0_1[15 : 8];
  assign zero_0_2 = tmp_zero_0_0_1[23 : 16];
  assign zero_0_3 = tmp_zero_0_0_1[31 : 24];
  assign zero_0_4 = tmp_zero_0_0_1[39 : 32];
  assign zero_0_5 = tmp_zero_0_0_1[47 : 40];
  assign zero_0_6 = tmp_zero_0_0_1[55 : 48];
  assign zero_0_7 = tmp_zero_0_0_1[63 : 56];
  assign zero_0_8 = tmp_zero_0_0_1[71 : 64];
  assign zero_0_9 = tmp_zero_0_0_1[79 : 72];
  assign zero_0_10 = tmp_zero_0_0_1[87 : 80];
  assign zero_0_11 = tmp_zero_0_0_1[95 : 88];
  assign zero_0_12 = tmp_zero_0_0_1[103 : 96];
  assign zero_0_13 = tmp_zero_0_0_1[111 : 104];
  assign zero_0_14 = tmp_zero_0_0_1[119 : 112];
  assign zero_0_15 = tmp_zero_0_0_1[127 : 120];
  assign tmp_zero_1_0 = tmp_zero_0_0[255 : 128];
  assign zero_1_0 = tmp_zero_1_0[7 : 0];
  assign zero_1_1 = tmp_zero_1_0[15 : 8];
  assign zero_1_2 = tmp_zero_1_0[23 : 16];
  assign zero_1_3 = tmp_zero_1_0[31 : 24];
  assign zero_1_4 = tmp_zero_1_0[39 : 32];
  assign zero_1_5 = tmp_zero_1_0[47 : 40];
  assign zero_1_6 = tmp_zero_1_0[55 : 48];
  assign zero_1_7 = tmp_zero_1_0[63 : 56];
  assign zero_1_8 = tmp_zero_1_0[71 : 64];
  assign zero_1_9 = tmp_zero_1_0[79 : 72];
  assign zero_1_10 = tmp_zero_1_0[87 : 80];
  assign zero_1_11 = tmp_zero_1_0[95 : 88];
  assign zero_1_12 = tmp_zero_1_0[103 : 96];
  assign zero_1_13 = tmp_zero_1_0[111 : 104];
  assign zero_1_14 = tmp_zero_1_0[119 : 112];
  assign zero_1_15 = tmp_zero_1_0[127 : 120];
  assign tmp_zero_2_0 = tmp_zero_0_0[383 : 256];
  assign zero_2_0 = tmp_zero_2_0[7 : 0];
  assign zero_2_1 = tmp_zero_2_0[15 : 8];
  assign zero_2_2 = tmp_zero_2_0[23 : 16];
  assign zero_2_3 = tmp_zero_2_0[31 : 24];
  assign zero_2_4 = tmp_zero_2_0[39 : 32];
  assign zero_2_5 = tmp_zero_2_0[47 : 40];
  assign zero_2_6 = tmp_zero_2_0[55 : 48];
  assign zero_2_7 = tmp_zero_2_0[63 : 56];
  assign zero_2_8 = tmp_zero_2_0[71 : 64];
  assign zero_2_9 = tmp_zero_2_0[79 : 72];
  assign zero_2_10 = tmp_zero_2_0[87 : 80];
  assign zero_2_11 = tmp_zero_2_0[95 : 88];
  assign zero_2_12 = tmp_zero_2_0[103 : 96];
  assign zero_2_13 = tmp_zero_2_0[111 : 104];
  assign zero_2_14 = tmp_zero_2_0[119 : 112];
  assign zero_2_15 = tmp_zero_2_0[127 : 120];
  assign videoInFire = (videoIn_valid && videoIn_ready);
  assign videoOutFire = (videoOut_valid && videoOut_ready);
  assign paddedFire = (padded_valid && padded_ready);
  assign when_PixelBufferSame_l46 = (videoInFire && videoIn_payload_endOfPack);
  always @(*) begin
    tmp_bridge_payload_endOfPack = 1'b0;
    if(when_PixelBufferSame_l48) begin
      tmp_bridge_payload_endOfPack = 1'b1;
    end
  end

  assign tmp_bridge_payload_endOfPack_1 = 1'b1;
  assign tmp_bridge_payload_endOfPack_2 = (tmp_bridge_payload_endOfPack_1 && tmp_bridge_payload_endOfPack);
  assign when_PixelBufferSame_l48 = (paddedFire && paddedCond);
  always @(*) begin
    tmp_padded_valid = videoIn_valid;
    if(paddedCond) begin
      tmp_padded_valid = 1'b1;
    end
  end

  always @(*) begin
    videoIn_ready = padded_ready;
    if(paddedCond) begin
      videoIn_ready = 1'b0;
    end
  end

  assign padded_valid = tmp_padded_valid;
  assign padded_payload_frame_line_pixel_0_0 = videoIn_payload_frame_line_pixel_0_0;
  assign padded_payload_frame_line_pixel_0_1 = videoIn_payload_frame_line_pixel_0_1;
  assign padded_payload_frame_line_pixel_0_2 = videoIn_payload_frame_line_pixel_0_2;
  assign padded_payload_frame_line_pixel_0_3 = videoIn_payload_frame_line_pixel_0_3;
  assign padded_payload_frame_line_pixel_0_4 = videoIn_payload_frame_line_pixel_0_4;
  assign padded_payload_frame_line_pixel_0_5 = videoIn_payload_frame_line_pixel_0_5;
  assign padded_payload_frame_line_pixel_0_6 = videoIn_payload_frame_line_pixel_0_6;
  assign padded_payload_frame_line_pixel_0_7 = videoIn_payload_frame_line_pixel_0_7;
  assign padded_payload_frame_line_pixel_0_8 = videoIn_payload_frame_line_pixel_0_8;
  assign padded_payload_frame_line_pixel_0_9 = videoIn_payload_frame_line_pixel_0_9;
  assign padded_payload_frame_line_pixel_0_10 = videoIn_payload_frame_line_pixel_0_10;
  assign padded_payload_frame_line_pixel_0_11 = videoIn_payload_frame_line_pixel_0_11;
  assign padded_payload_frame_line_pixel_0_12 = videoIn_payload_frame_line_pixel_0_12;
  assign padded_payload_frame_line_pixel_0_13 = videoIn_payload_frame_line_pixel_0_13;
  assign padded_payload_frame_line_pixel_0_14 = videoIn_payload_frame_line_pixel_0_14;
  assign padded_payload_frame_line_pixel_0_15 = videoIn_payload_frame_line_pixel_0_15;
  assign padded_payload_frame_line_pixel_1_0 = videoIn_payload_frame_line_pixel_1_0;
  assign padded_payload_frame_line_pixel_1_1 = videoIn_payload_frame_line_pixel_1_1;
  assign padded_payload_frame_line_pixel_1_2 = videoIn_payload_frame_line_pixel_1_2;
  assign padded_payload_frame_line_pixel_1_3 = videoIn_payload_frame_line_pixel_1_3;
  assign padded_payload_frame_line_pixel_1_4 = videoIn_payload_frame_line_pixel_1_4;
  assign padded_payload_frame_line_pixel_1_5 = videoIn_payload_frame_line_pixel_1_5;
  assign padded_payload_frame_line_pixel_1_6 = videoIn_payload_frame_line_pixel_1_6;
  assign padded_payload_frame_line_pixel_1_7 = videoIn_payload_frame_line_pixel_1_7;
  assign padded_payload_frame_line_pixel_1_8 = videoIn_payload_frame_line_pixel_1_8;
  assign padded_payload_frame_line_pixel_1_9 = videoIn_payload_frame_line_pixel_1_9;
  assign padded_payload_frame_line_pixel_1_10 = videoIn_payload_frame_line_pixel_1_10;
  assign padded_payload_frame_line_pixel_1_11 = videoIn_payload_frame_line_pixel_1_11;
  assign padded_payload_frame_line_pixel_1_12 = videoIn_payload_frame_line_pixel_1_12;
  assign padded_payload_frame_line_pixel_1_13 = videoIn_payload_frame_line_pixel_1_13;
  assign padded_payload_frame_line_pixel_1_14 = videoIn_payload_frame_line_pixel_1_14;
  assign padded_payload_frame_line_pixel_1_15 = videoIn_payload_frame_line_pixel_1_15;
  assign padded_payload_frame_line_pixel_2_0 = videoIn_payload_frame_line_pixel_2_0;
  assign padded_payload_frame_line_pixel_2_1 = videoIn_payload_frame_line_pixel_2_1;
  assign padded_payload_frame_line_pixel_2_2 = videoIn_payload_frame_line_pixel_2_2;
  assign padded_payload_frame_line_pixel_2_3 = videoIn_payload_frame_line_pixel_2_3;
  assign padded_payload_frame_line_pixel_2_4 = videoIn_payload_frame_line_pixel_2_4;
  assign padded_payload_frame_line_pixel_2_5 = videoIn_payload_frame_line_pixel_2_5;
  assign padded_payload_frame_line_pixel_2_6 = videoIn_payload_frame_line_pixel_2_6;
  assign padded_payload_frame_line_pixel_2_7 = videoIn_payload_frame_line_pixel_2_7;
  assign padded_payload_frame_line_pixel_2_8 = videoIn_payload_frame_line_pixel_2_8;
  assign padded_payload_frame_line_pixel_2_9 = videoIn_payload_frame_line_pixel_2_9;
  assign padded_payload_frame_line_pixel_2_10 = videoIn_payload_frame_line_pixel_2_10;
  assign padded_payload_frame_line_pixel_2_11 = videoIn_payload_frame_line_pixel_2_11;
  assign padded_payload_frame_line_pixel_2_12 = videoIn_payload_frame_line_pixel_2_12;
  assign padded_payload_frame_line_pixel_2_13 = videoIn_payload_frame_line_pixel_2_13;
  assign padded_payload_frame_line_pixel_2_14 = videoIn_payload_frame_line_pixel_2_14;
  assign padded_payload_frame_line_pixel_2_15 = videoIn_payload_frame_line_pixel_2_15;
  assign padded_payload_frame_line_endOfLine = videoIn_payload_frame_line_endOfLine;
  assign padded_payload_frame_endOfFrame = videoIn_payload_frame_endOfFrame;
  assign padded_payload_endOfPack = videoIn_payload_endOfPack;
  assign bridgeFire = (bridge_valid && bridge_ready);
  assign bridge_valid = padded_valid;
  assign padded_ready = bridge_ready;
  assign cntPrevStable = (cntPrev == 2'b01);
  assign cntPostStable = (cntPost == 2'b01);
  assign cntPrevEqualVec_0 = ((2'b00 <= cntPrev) && (cntPrev < 2'b01));
  assign cntPostEqualVec_0 = (cntPost <= 2'b00);
  assign when_PixelBufferSame_l74 = (videoInFire && videoIn_payload_frame_line_endOfLine);
  assign when_PixelBufferSame_l75 = (videoOutFire && videoOut_payload_frame_line_endOfLine);
  assign when_PixelBufferSame_l76 = (videoOutFire && (! cntPrevStable));
  assign when_PixelBufferSame_l77 = (videoOutFire && (! cntPostStable));
  assign tmp_pixelVec_0_0_0 = {{{videoIn_payload_frame_line_pixel_2_15,{videoIn_payload_frame_line_pixel_2_14,{videoIn_payload_frame_line_pixel_2_13,{videoIn_payload_frame_line_pixel_2_12,{tmp_tmp_pixelVec_0_0_0,tmp_tmp_pixelVec_0_0_0_1}}}}},{{videoIn_payload_frame_line_pixel_1_15,{videoIn_payload_frame_line_pixel_1_14,{videoIn_payload_frame_line_pixel_1_13,{tmp_tmp_pixelVec_0_0_0_4,tmp_tmp_pixelVec_0_0_0_5}}}},{videoIn_payload_frame_line_pixel_0_15,{videoIn_payload_frame_line_pixel_0_14,{videoIn_payload_frame_line_pixel_0_13,{tmp_tmp_pixelVec_0_0_0_8,tmp_tmp_pixelVec_0_0_0_9}}}}}},pixelBuffer};
  assign tmp_pixelVec_0_0_0_1 = tmp_pixelVec_0_0_0[383 : 0];
  assign tmp_pixelVec_0_0_0_2 = tmp_pixelVec_0_0_0_1[127 : 0];
  assign pixelVec_0_0_0 = tmp_pixelVec_0_0_0_2[7 : 0];
  assign pixelVec_0_0_1 = tmp_pixelVec_0_0_0_2[15 : 8];
  assign pixelVec_0_0_2 = tmp_pixelVec_0_0_0_2[23 : 16];
  assign pixelVec_0_0_3 = tmp_pixelVec_0_0_0_2[31 : 24];
  assign pixelVec_0_0_4 = tmp_pixelVec_0_0_0_2[39 : 32];
  assign pixelVec_0_0_5 = tmp_pixelVec_0_0_0_2[47 : 40];
  assign pixelVec_0_0_6 = tmp_pixelVec_0_0_0_2[55 : 48];
  assign pixelVec_0_0_7 = tmp_pixelVec_0_0_0_2[63 : 56];
  assign pixelVec_0_0_8 = tmp_pixelVec_0_0_0_2[71 : 64];
  assign pixelVec_0_0_9 = tmp_pixelVec_0_0_0_2[79 : 72];
  assign pixelVec_0_0_10 = tmp_pixelVec_0_0_0_2[87 : 80];
  assign pixelVec_0_0_11 = tmp_pixelVec_0_0_0_2[95 : 88];
  assign pixelVec_0_0_12 = tmp_pixelVec_0_0_0_2[103 : 96];
  assign pixelVec_0_0_13 = tmp_pixelVec_0_0_0_2[111 : 104];
  assign pixelVec_0_0_14 = tmp_pixelVec_0_0_0_2[119 : 112];
  assign pixelVec_0_0_15 = tmp_pixelVec_0_0_0_2[127 : 120];
  assign tmp_pixelVec_0_1_0 = tmp_pixelVec_0_0_0_1[255 : 128];
  assign pixelVec_0_1_0 = tmp_pixelVec_0_1_0[7 : 0];
  assign pixelVec_0_1_1 = tmp_pixelVec_0_1_0[15 : 8];
  assign pixelVec_0_1_2 = tmp_pixelVec_0_1_0[23 : 16];
  assign pixelVec_0_1_3 = tmp_pixelVec_0_1_0[31 : 24];
  assign pixelVec_0_1_4 = tmp_pixelVec_0_1_0[39 : 32];
  assign pixelVec_0_1_5 = tmp_pixelVec_0_1_0[47 : 40];
  assign pixelVec_0_1_6 = tmp_pixelVec_0_1_0[55 : 48];
  assign pixelVec_0_1_7 = tmp_pixelVec_0_1_0[63 : 56];
  assign pixelVec_0_1_8 = tmp_pixelVec_0_1_0[71 : 64];
  assign pixelVec_0_1_9 = tmp_pixelVec_0_1_0[79 : 72];
  assign pixelVec_0_1_10 = tmp_pixelVec_0_1_0[87 : 80];
  assign pixelVec_0_1_11 = tmp_pixelVec_0_1_0[95 : 88];
  assign pixelVec_0_1_12 = tmp_pixelVec_0_1_0[103 : 96];
  assign pixelVec_0_1_13 = tmp_pixelVec_0_1_0[111 : 104];
  assign pixelVec_0_1_14 = tmp_pixelVec_0_1_0[119 : 112];
  assign pixelVec_0_1_15 = tmp_pixelVec_0_1_0[127 : 120];
  assign tmp_pixelVec_0_2_0 = tmp_pixelVec_0_0_0_1[383 : 256];
  assign pixelVec_0_2_0 = tmp_pixelVec_0_2_0[7 : 0];
  assign pixelVec_0_2_1 = tmp_pixelVec_0_2_0[15 : 8];
  assign pixelVec_0_2_2 = tmp_pixelVec_0_2_0[23 : 16];
  assign pixelVec_0_2_3 = tmp_pixelVec_0_2_0[31 : 24];
  assign pixelVec_0_2_4 = tmp_pixelVec_0_2_0[39 : 32];
  assign pixelVec_0_2_5 = tmp_pixelVec_0_2_0[47 : 40];
  assign pixelVec_0_2_6 = tmp_pixelVec_0_2_0[55 : 48];
  assign pixelVec_0_2_7 = tmp_pixelVec_0_2_0[63 : 56];
  assign pixelVec_0_2_8 = tmp_pixelVec_0_2_0[71 : 64];
  assign pixelVec_0_2_9 = tmp_pixelVec_0_2_0[79 : 72];
  assign pixelVec_0_2_10 = tmp_pixelVec_0_2_0[87 : 80];
  assign pixelVec_0_2_11 = tmp_pixelVec_0_2_0[95 : 88];
  assign pixelVec_0_2_12 = tmp_pixelVec_0_2_0[103 : 96];
  assign pixelVec_0_2_13 = tmp_pixelVec_0_2_0[111 : 104];
  assign pixelVec_0_2_14 = tmp_pixelVec_0_2_0[119 : 112];
  assign pixelVec_0_2_15 = tmp_pixelVec_0_2_0[127 : 120];
  assign tmp_pixelVec_1_0_0 = tmp_pixelVec_0_0_0[767 : 384];
  assign tmp_pixelVec_1_0_0_1 = tmp_pixelVec_1_0_0[127 : 0];
  assign pixelVec_1_0_0 = tmp_pixelVec_1_0_0_1[7 : 0];
  assign pixelVec_1_0_1 = tmp_pixelVec_1_0_0_1[15 : 8];
  assign pixelVec_1_0_2 = tmp_pixelVec_1_0_0_1[23 : 16];
  assign pixelVec_1_0_3 = tmp_pixelVec_1_0_0_1[31 : 24];
  assign pixelVec_1_0_4 = tmp_pixelVec_1_0_0_1[39 : 32];
  assign pixelVec_1_0_5 = tmp_pixelVec_1_0_0_1[47 : 40];
  assign pixelVec_1_0_6 = tmp_pixelVec_1_0_0_1[55 : 48];
  assign pixelVec_1_0_7 = tmp_pixelVec_1_0_0_1[63 : 56];
  assign pixelVec_1_0_8 = tmp_pixelVec_1_0_0_1[71 : 64];
  assign pixelVec_1_0_9 = tmp_pixelVec_1_0_0_1[79 : 72];
  assign pixelVec_1_0_10 = tmp_pixelVec_1_0_0_1[87 : 80];
  assign pixelVec_1_0_11 = tmp_pixelVec_1_0_0_1[95 : 88];
  assign pixelVec_1_0_12 = tmp_pixelVec_1_0_0_1[103 : 96];
  assign pixelVec_1_0_13 = tmp_pixelVec_1_0_0_1[111 : 104];
  assign pixelVec_1_0_14 = tmp_pixelVec_1_0_0_1[119 : 112];
  assign pixelVec_1_0_15 = tmp_pixelVec_1_0_0_1[127 : 120];
  assign tmp_pixelVec_1_1_0 = tmp_pixelVec_1_0_0[255 : 128];
  assign pixelVec_1_1_0 = tmp_pixelVec_1_1_0[7 : 0];
  assign pixelVec_1_1_1 = tmp_pixelVec_1_1_0[15 : 8];
  assign pixelVec_1_1_2 = tmp_pixelVec_1_1_0[23 : 16];
  assign pixelVec_1_1_3 = tmp_pixelVec_1_1_0[31 : 24];
  assign pixelVec_1_1_4 = tmp_pixelVec_1_1_0[39 : 32];
  assign pixelVec_1_1_5 = tmp_pixelVec_1_1_0[47 : 40];
  assign pixelVec_1_1_6 = tmp_pixelVec_1_1_0[55 : 48];
  assign pixelVec_1_1_7 = tmp_pixelVec_1_1_0[63 : 56];
  assign pixelVec_1_1_8 = tmp_pixelVec_1_1_0[71 : 64];
  assign pixelVec_1_1_9 = tmp_pixelVec_1_1_0[79 : 72];
  assign pixelVec_1_1_10 = tmp_pixelVec_1_1_0[87 : 80];
  assign pixelVec_1_1_11 = tmp_pixelVec_1_1_0[95 : 88];
  assign pixelVec_1_1_12 = tmp_pixelVec_1_1_0[103 : 96];
  assign pixelVec_1_1_13 = tmp_pixelVec_1_1_0[111 : 104];
  assign pixelVec_1_1_14 = tmp_pixelVec_1_1_0[119 : 112];
  assign pixelVec_1_1_15 = tmp_pixelVec_1_1_0[127 : 120];
  assign tmp_pixelVec_1_2_0 = tmp_pixelVec_1_0_0[383 : 256];
  assign pixelVec_1_2_0 = tmp_pixelVec_1_2_0[7 : 0];
  assign pixelVec_1_2_1 = tmp_pixelVec_1_2_0[15 : 8];
  assign pixelVec_1_2_2 = tmp_pixelVec_1_2_0[23 : 16];
  assign pixelVec_1_2_3 = tmp_pixelVec_1_2_0[31 : 24];
  assign pixelVec_1_2_4 = tmp_pixelVec_1_2_0[39 : 32];
  assign pixelVec_1_2_5 = tmp_pixelVec_1_2_0[47 : 40];
  assign pixelVec_1_2_6 = tmp_pixelVec_1_2_0[55 : 48];
  assign pixelVec_1_2_7 = tmp_pixelVec_1_2_0[63 : 56];
  assign pixelVec_1_2_8 = tmp_pixelVec_1_2_0[71 : 64];
  assign pixelVec_1_2_9 = tmp_pixelVec_1_2_0[79 : 72];
  assign pixelVec_1_2_10 = tmp_pixelVec_1_2_0[87 : 80];
  assign pixelVec_1_2_11 = tmp_pixelVec_1_2_0[95 : 88];
  assign pixelVec_1_2_12 = tmp_pixelVec_1_2_0[103 : 96];
  assign pixelVec_1_2_13 = tmp_pixelVec_1_2_0[111 : 104];
  assign pixelVec_1_2_14 = tmp_pixelVec_1_2_0[119 : 112];
  assign pixelVec_1_2_15 = tmp_pixelVec_1_2_0[127 : 120];
  assign tmp_pixelVec_2_0_0 = tmp_pixelVec_0_0_0[1151 : 768];
  assign tmp_pixelVec_2_0_0_1 = tmp_pixelVec_2_0_0[127 : 0];
  assign pixelVec_2_0_0 = tmp_pixelVec_2_0_0_1[7 : 0];
  assign pixelVec_2_0_1 = tmp_pixelVec_2_0_0_1[15 : 8];
  assign pixelVec_2_0_2 = tmp_pixelVec_2_0_0_1[23 : 16];
  assign pixelVec_2_0_3 = tmp_pixelVec_2_0_0_1[31 : 24];
  assign pixelVec_2_0_4 = tmp_pixelVec_2_0_0_1[39 : 32];
  assign pixelVec_2_0_5 = tmp_pixelVec_2_0_0_1[47 : 40];
  assign pixelVec_2_0_6 = tmp_pixelVec_2_0_0_1[55 : 48];
  assign pixelVec_2_0_7 = tmp_pixelVec_2_0_0_1[63 : 56];
  assign pixelVec_2_0_8 = tmp_pixelVec_2_0_0_1[71 : 64];
  assign pixelVec_2_0_9 = tmp_pixelVec_2_0_0_1[79 : 72];
  assign pixelVec_2_0_10 = tmp_pixelVec_2_0_0_1[87 : 80];
  assign pixelVec_2_0_11 = tmp_pixelVec_2_0_0_1[95 : 88];
  assign pixelVec_2_0_12 = tmp_pixelVec_2_0_0_1[103 : 96];
  assign pixelVec_2_0_13 = tmp_pixelVec_2_0_0_1[111 : 104];
  assign pixelVec_2_0_14 = tmp_pixelVec_2_0_0_1[119 : 112];
  assign pixelVec_2_0_15 = tmp_pixelVec_2_0_0_1[127 : 120];
  assign tmp_pixelVec_2_1_0 = tmp_pixelVec_2_0_0[255 : 128];
  assign pixelVec_2_1_0 = tmp_pixelVec_2_1_0[7 : 0];
  assign pixelVec_2_1_1 = tmp_pixelVec_2_1_0[15 : 8];
  assign pixelVec_2_1_2 = tmp_pixelVec_2_1_0[23 : 16];
  assign pixelVec_2_1_3 = tmp_pixelVec_2_1_0[31 : 24];
  assign pixelVec_2_1_4 = tmp_pixelVec_2_1_0[39 : 32];
  assign pixelVec_2_1_5 = tmp_pixelVec_2_1_0[47 : 40];
  assign pixelVec_2_1_6 = tmp_pixelVec_2_1_0[55 : 48];
  assign pixelVec_2_1_7 = tmp_pixelVec_2_1_0[63 : 56];
  assign pixelVec_2_1_8 = tmp_pixelVec_2_1_0[71 : 64];
  assign pixelVec_2_1_9 = tmp_pixelVec_2_1_0[79 : 72];
  assign pixelVec_2_1_10 = tmp_pixelVec_2_1_0[87 : 80];
  assign pixelVec_2_1_11 = tmp_pixelVec_2_1_0[95 : 88];
  assign pixelVec_2_1_12 = tmp_pixelVec_2_1_0[103 : 96];
  assign pixelVec_2_1_13 = tmp_pixelVec_2_1_0[111 : 104];
  assign pixelVec_2_1_14 = tmp_pixelVec_2_1_0[119 : 112];
  assign pixelVec_2_1_15 = tmp_pixelVec_2_1_0[127 : 120];
  assign tmp_pixelVec_2_2_0 = tmp_pixelVec_2_0_0[383 : 256];
  assign pixelVec_2_2_0 = tmp_pixelVec_2_2_0[7 : 0];
  assign pixelVec_2_2_1 = tmp_pixelVec_2_2_0[15 : 8];
  assign pixelVec_2_2_2 = tmp_pixelVec_2_2_0[23 : 16];
  assign pixelVec_2_2_3 = tmp_pixelVec_2_2_0[31 : 24];
  assign pixelVec_2_2_4 = tmp_pixelVec_2_2_0[39 : 32];
  assign pixelVec_2_2_5 = tmp_pixelVec_2_2_0[47 : 40];
  assign pixelVec_2_2_6 = tmp_pixelVec_2_2_0[55 : 48];
  assign pixelVec_2_2_7 = tmp_pixelVec_2_2_0[63 : 56];
  assign pixelVec_2_2_8 = tmp_pixelVec_2_2_0[71 : 64];
  assign pixelVec_2_2_9 = tmp_pixelVec_2_2_0[79 : 72];
  assign pixelVec_2_2_10 = tmp_pixelVec_2_2_0[87 : 80];
  assign pixelVec_2_2_11 = tmp_pixelVec_2_2_0[95 : 88];
  assign pixelVec_2_2_12 = tmp_pixelVec_2_2_0[103 : 96];
  assign pixelVec_2_2_13 = tmp_pixelVec_2_2_0[111 : 104];
  assign pixelVec_2_2_14 = tmp_pixelVec_2_2_0[119 : 112];
  assign pixelVec_2_2_15 = tmp_pixelVec_2_2_0[127 : 120];
  assign up_0_0_0 = (cntPostEqualVec_0 ? zero_0_0 : pixelVec_0_0_0);
  assign up_0_0_1 = (cntPostEqualVec_0 ? zero_0_1 : pixelVec_0_0_1);
  assign up_0_0_2 = (cntPostEqualVec_0 ? zero_0_2 : pixelVec_0_0_2);
  assign up_0_0_3 = (cntPostEqualVec_0 ? zero_0_3 : pixelVec_0_0_3);
  assign up_0_0_4 = (cntPostEqualVec_0 ? zero_0_4 : pixelVec_0_0_4);
  assign up_0_0_5 = (cntPostEqualVec_0 ? zero_0_5 : pixelVec_0_0_5);
  assign up_0_0_6 = (cntPostEqualVec_0 ? zero_0_6 : pixelVec_0_0_6);
  assign up_0_0_7 = (cntPostEqualVec_0 ? zero_0_7 : pixelVec_0_0_7);
  assign up_0_0_8 = (cntPostEqualVec_0 ? zero_0_8 : pixelVec_0_0_8);
  assign up_0_0_9 = (cntPostEqualVec_0 ? zero_0_9 : pixelVec_0_0_9);
  assign up_0_0_10 = (cntPostEqualVec_0 ? zero_0_10 : pixelVec_0_0_10);
  assign up_0_0_11 = (cntPostEqualVec_0 ? zero_0_11 : pixelVec_0_0_11);
  assign up_0_0_12 = (cntPostEqualVec_0 ? zero_0_12 : pixelVec_0_0_12);
  assign up_0_0_13 = (cntPostEqualVec_0 ? zero_0_13 : pixelVec_0_0_13);
  assign up_0_0_14 = (cntPostEqualVec_0 ? zero_0_14 : pixelVec_0_0_14);
  assign up_0_0_15 = (cntPostEqualVec_0 ? zero_0_15 : pixelVec_0_0_15);
  assign up_0_1_0 = (cntPostEqualVec_0 ? zero_1_0 : pixelVec_0_1_0);
  assign up_0_1_1 = (cntPostEqualVec_0 ? zero_1_1 : pixelVec_0_1_1);
  assign up_0_1_2 = (cntPostEqualVec_0 ? zero_1_2 : pixelVec_0_1_2);
  assign up_0_1_3 = (cntPostEqualVec_0 ? zero_1_3 : pixelVec_0_1_3);
  assign up_0_1_4 = (cntPostEqualVec_0 ? zero_1_4 : pixelVec_0_1_4);
  assign up_0_1_5 = (cntPostEqualVec_0 ? zero_1_5 : pixelVec_0_1_5);
  assign up_0_1_6 = (cntPostEqualVec_0 ? zero_1_6 : pixelVec_0_1_6);
  assign up_0_1_7 = (cntPostEqualVec_0 ? zero_1_7 : pixelVec_0_1_7);
  assign up_0_1_8 = (cntPostEqualVec_0 ? zero_1_8 : pixelVec_0_1_8);
  assign up_0_1_9 = (cntPostEqualVec_0 ? zero_1_9 : pixelVec_0_1_9);
  assign up_0_1_10 = (cntPostEqualVec_0 ? zero_1_10 : pixelVec_0_1_10);
  assign up_0_1_11 = (cntPostEqualVec_0 ? zero_1_11 : pixelVec_0_1_11);
  assign up_0_1_12 = (cntPostEqualVec_0 ? zero_1_12 : pixelVec_0_1_12);
  assign up_0_1_13 = (cntPostEqualVec_0 ? zero_1_13 : pixelVec_0_1_13);
  assign up_0_1_14 = (cntPostEqualVec_0 ? zero_1_14 : pixelVec_0_1_14);
  assign up_0_1_15 = (cntPostEqualVec_0 ? zero_1_15 : pixelVec_0_1_15);
  assign up_0_2_0 = (cntPostEqualVec_0 ? zero_2_0 : pixelVec_0_2_0);
  assign up_0_2_1 = (cntPostEqualVec_0 ? zero_2_1 : pixelVec_0_2_1);
  assign up_0_2_2 = (cntPostEqualVec_0 ? zero_2_2 : pixelVec_0_2_2);
  assign up_0_2_3 = (cntPostEqualVec_0 ? zero_2_3 : pixelVec_0_2_3);
  assign up_0_2_4 = (cntPostEqualVec_0 ? zero_2_4 : pixelVec_0_2_4);
  assign up_0_2_5 = (cntPostEqualVec_0 ? zero_2_5 : pixelVec_0_2_5);
  assign up_0_2_6 = (cntPostEqualVec_0 ? zero_2_6 : pixelVec_0_2_6);
  assign up_0_2_7 = (cntPostEqualVec_0 ? zero_2_7 : pixelVec_0_2_7);
  assign up_0_2_8 = (cntPostEqualVec_0 ? zero_2_8 : pixelVec_0_2_8);
  assign up_0_2_9 = (cntPostEqualVec_0 ? zero_2_9 : pixelVec_0_2_9);
  assign up_0_2_10 = (cntPostEqualVec_0 ? zero_2_10 : pixelVec_0_2_10);
  assign up_0_2_11 = (cntPostEqualVec_0 ? zero_2_11 : pixelVec_0_2_11);
  assign up_0_2_12 = (cntPostEqualVec_0 ? zero_2_12 : pixelVec_0_2_12);
  assign up_0_2_13 = (cntPostEqualVec_0 ? zero_2_13 : pixelVec_0_2_13);
  assign up_0_2_14 = (cntPostEqualVec_0 ? zero_2_14 : pixelVec_0_2_14);
  assign up_0_2_15 = (cntPostEqualVec_0 ? zero_2_15 : pixelVec_0_2_15);
  assign down_0_0_0 = (cntPrevEqualVec_0 ? zero_0_0 : pixelVec_2_0_0);
  assign down_0_0_1 = (cntPrevEqualVec_0 ? zero_0_1 : pixelVec_2_0_1);
  assign down_0_0_2 = (cntPrevEqualVec_0 ? zero_0_2 : pixelVec_2_0_2);
  assign down_0_0_3 = (cntPrevEqualVec_0 ? zero_0_3 : pixelVec_2_0_3);
  assign down_0_0_4 = (cntPrevEqualVec_0 ? zero_0_4 : pixelVec_2_0_4);
  assign down_0_0_5 = (cntPrevEqualVec_0 ? zero_0_5 : pixelVec_2_0_5);
  assign down_0_0_6 = (cntPrevEqualVec_0 ? zero_0_6 : pixelVec_2_0_6);
  assign down_0_0_7 = (cntPrevEqualVec_0 ? zero_0_7 : pixelVec_2_0_7);
  assign down_0_0_8 = (cntPrevEqualVec_0 ? zero_0_8 : pixelVec_2_0_8);
  assign down_0_0_9 = (cntPrevEqualVec_0 ? zero_0_9 : pixelVec_2_0_9);
  assign down_0_0_10 = (cntPrevEqualVec_0 ? zero_0_10 : pixelVec_2_0_10);
  assign down_0_0_11 = (cntPrevEqualVec_0 ? zero_0_11 : pixelVec_2_0_11);
  assign down_0_0_12 = (cntPrevEqualVec_0 ? zero_0_12 : pixelVec_2_0_12);
  assign down_0_0_13 = (cntPrevEqualVec_0 ? zero_0_13 : pixelVec_2_0_13);
  assign down_0_0_14 = (cntPrevEqualVec_0 ? zero_0_14 : pixelVec_2_0_14);
  assign down_0_0_15 = (cntPrevEqualVec_0 ? zero_0_15 : pixelVec_2_0_15);
  assign down_0_1_0 = (cntPrevEqualVec_0 ? zero_1_0 : pixelVec_2_1_0);
  assign down_0_1_1 = (cntPrevEqualVec_0 ? zero_1_1 : pixelVec_2_1_1);
  assign down_0_1_2 = (cntPrevEqualVec_0 ? zero_1_2 : pixelVec_2_1_2);
  assign down_0_1_3 = (cntPrevEqualVec_0 ? zero_1_3 : pixelVec_2_1_3);
  assign down_0_1_4 = (cntPrevEqualVec_0 ? zero_1_4 : pixelVec_2_1_4);
  assign down_0_1_5 = (cntPrevEqualVec_0 ? zero_1_5 : pixelVec_2_1_5);
  assign down_0_1_6 = (cntPrevEqualVec_0 ? zero_1_6 : pixelVec_2_1_6);
  assign down_0_1_7 = (cntPrevEqualVec_0 ? zero_1_7 : pixelVec_2_1_7);
  assign down_0_1_8 = (cntPrevEqualVec_0 ? zero_1_8 : pixelVec_2_1_8);
  assign down_0_1_9 = (cntPrevEqualVec_0 ? zero_1_9 : pixelVec_2_1_9);
  assign down_0_1_10 = (cntPrevEqualVec_0 ? zero_1_10 : pixelVec_2_1_10);
  assign down_0_1_11 = (cntPrevEqualVec_0 ? zero_1_11 : pixelVec_2_1_11);
  assign down_0_1_12 = (cntPrevEqualVec_0 ? zero_1_12 : pixelVec_2_1_12);
  assign down_0_1_13 = (cntPrevEqualVec_0 ? zero_1_13 : pixelVec_2_1_13);
  assign down_0_1_14 = (cntPrevEqualVec_0 ? zero_1_14 : pixelVec_2_1_14);
  assign down_0_1_15 = (cntPrevEqualVec_0 ? zero_1_15 : pixelVec_2_1_15);
  assign down_0_2_0 = (cntPrevEqualVec_0 ? zero_2_0 : pixelVec_2_2_0);
  assign down_0_2_1 = (cntPrevEqualVec_0 ? zero_2_1 : pixelVec_2_2_1);
  assign down_0_2_2 = (cntPrevEqualVec_0 ? zero_2_2 : pixelVec_2_2_2);
  assign down_0_2_3 = (cntPrevEqualVec_0 ? zero_2_3 : pixelVec_2_2_3);
  assign down_0_2_4 = (cntPrevEqualVec_0 ? zero_2_4 : pixelVec_2_2_4);
  assign down_0_2_5 = (cntPrevEqualVec_0 ? zero_2_5 : pixelVec_2_2_5);
  assign down_0_2_6 = (cntPrevEqualVec_0 ? zero_2_6 : pixelVec_2_2_6);
  assign down_0_2_7 = (cntPrevEqualVec_0 ? zero_2_7 : pixelVec_2_2_7);
  assign down_0_2_8 = (cntPrevEqualVec_0 ? zero_2_8 : pixelVec_2_2_8);
  assign down_0_2_9 = (cntPrevEqualVec_0 ? zero_2_9 : pixelVec_2_2_9);
  assign down_0_2_10 = (cntPrevEqualVec_0 ? zero_2_10 : pixelVec_2_2_10);
  assign down_0_2_11 = (cntPrevEqualVec_0 ? zero_2_11 : pixelVec_2_2_11);
  assign down_0_2_12 = (cntPrevEqualVec_0 ? zero_2_12 : pixelVec_2_2_12);
  assign down_0_2_13 = (cntPrevEqualVec_0 ? zero_2_13 : pixelVec_2_2_13);
  assign down_0_2_14 = (cntPrevEqualVec_0 ? zero_2_14 : pixelVec_2_2_14);
  assign down_0_2_15 = (cntPrevEqualVec_0 ? zero_2_15 : pixelVec_2_2_15);
  assign bridge_payload_endOfPack = tmp_bridge_payload_endOfPack_2;
  assign bridge_payload_frame_endOfFrame = padded_payload_frame_endOfFrame_delay_1;
  assign bridge_payload_frame_line_endOfLine = padded_payload_frame_line_endOfLine_delay_1;
  assign bridge_payload_frame_line_pixel_0_0_0 = up_0_0_0;
  assign bridge_payload_frame_line_pixel_0_0_1 = up_0_0_1;
  assign bridge_payload_frame_line_pixel_0_0_2 = up_0_0_2;
  assign bridge_payload_frame_line_pixel_0_0_3 = up_0_0_3;
  assign bridge_payload_frame_line_pixel_0_0_4 = up_0_0_4;
  assign bridge_payload_frame_line_pixel_0_0_5 = up_0_0_5;
  assign bridge_payload_frame_line_pixel_0_0_6 = up_0_0_6;
  assign bridge_payload_frame_line_pixel_0_0_7 = up_0_0_7;
  assign bridge_payload_frame_line_pixel_0_0_8 = up_0_0_8;
  assign bridge_payload_frame_line_pixel_0_0_9 = up_0_0_9;
  assign bridge_payload_frame_line_pixel_0_0_10 = up_0_0_10;
  assign bridge_payload_frame_line_pixel_0_0_11 = up_0_0_11;
  assign bridge_payload_frame_line_pixel_0_0_12 = up_0_0_12;
  assign bridge_payload_frame_line_pixel_0_0_13 = up_0_0_13;
  assign bridge_payload_frame_line_pixel_0_0_14 = up_0_0_14;
  assign bridge_payload_frame_line_pixel_0_0_15 = up_0_0_15;
  assign bridge_payload_frame_line_pixel_0_1_0 = up_0_1_0;
  assign bridge_payload_frame_line_pixel_0_1_1 = up_0_1_1;
  assign bridge_payload_frame_line_pixel_0_1_2 = up_0_1_2;
  assign bridge_payload_frame_line_pixel_0_1_3 = up_0_1_3;
  assign bridge_payload_frame_line_pixel_0_1_4 = up_0_1_4;
  assign bridge_payload_frame_line_pixel_0_1_5 = up_0_1_5;
  assign bridge_payload_frame_line_pixel_0_1_6 = up_0_1_6;
  assign bridge_payload_frame_line_pixel_0_1_7 = up_0_1_7;
  assign bridge_payload_frame_line_pixel_0_1_8 = up_0_1_8;
  assign bridge_payload_frame_line_pixel_0_1_9 = up_0_1_9;
  assign bridge_payload_frame_line_pixel_0_1_10 = up_0_1_10;
  assign bridge_payload_frame_line_pixel_0_1_11 = up_0_1_11;
  assign bridge_payload_frame_line_pixel_0_1_12 = up_0_1_12;
  assign bridge_payload_frame_line_pixel_0_1_13 = up_0_1_13;
  assign bridge_payload_frame_line_pixel_0_1_14 = up_0_1_14;
  assign bridge_payload_frame_line_pixel_0_1_15 = up_0_1_15;
  assign bridge_payload_frame_line_pixel_0_2_0 = up_0_2_0;
  assign bridge_payload_frame_line_pixel_0_2_1 = up_0_2_1;
  assign bridge_payload_frame_line_pixel_0_2_2 = up_0_2_2;
  assign bridge_payload_frame_line_pixel_0_2_3 = up_0_2_3;
  assign bridge_payload_frame_line_pixel_0_2_4 = up_0_2_4;
  assign bridge_payload_frame_line_pixel_0_2_5 = up_0_2_5;
  assign bridge_payload_frame_line_pixel_0_2_6 = up_0_2_6;
  assign bridge_payload_frame_line_pixel_0_2_7 = up_0_2_7;
  assign bridge_payload_frame_line_pixel_0_2_8 = up_0_2_8;
  assign bridge_payload_frame_line_pixel_0_2_9 = up_0_2_9;
  assign bridge_payload_frame_line_pixel_0_2_10 = up_0_2_10;
  assign bridge_payload_frame_line_pixel_0_2_11 = up_0_2_11;
  assign bridge_payload_frame_line_pixel_0_2_12 = up_0_2_12;
  assign bridge_payload_frame_line_pixel_0_2_13 = up_0_2_13;
  assign bridge_payload_frame_line_pixel_0_2_14 = up_0_2_14;
  assign bridge_payload_frame_line_pixel_0_2_15 = up_0_2_15;
  assign bridge_payload_frame_line_pixel_1_0_0 = pixelVec_1_0_0;
  assign bridge_payload_frame_line_pixel_1_0_1 = pixelVec_1_0_1;
  assign bridge_payload_frame_line_pixel_1_0_2 = pixelVec_1_0_2;
  assign bridge_payload_frame_line_pixel_1_0_3 = pixelVec_1_0_3;
  assign bridge_payload_frame_line_pixel_1_0_4 = pixelVec_1_0_4;
  assign bridge_payload_frame_line_pixel_1_0_5 = pixelVec_1_0_5;
  assign bridge_payload_frame_line_pixel_1_0_6 = pixelVec_1_0_6;
  assign bridge_payload_frame_line_pixel_1_0_7 = pixelVec_1_0_7;
  assign bridge_payload_frame_line_pixel_1_0_8 = pixelVec_1_0_8;
  assign bridge_payload_frame_line_pixel_1_0_9 = pixelVec_1_0_9;
  assign bridge_payload_frame_line_pixel_1_0_10 = pixelVec_1_0_10;
  assign bridge_payload_frame_line_pixel_1_0_11 = pixelVec_1_0_11;
  assign bridge_payload_frame_line_pixel_1_0_12 = pixelVec_1_0_12;
  assign bridge_payload_frame_line_pixel_1_0_13 = pixelVec_1_0_13;
  assign bridge_payload_frame_line_pixel_1_0_14 = pixelVec_1_0_14;
  assign bridge_payload_frame_line_pixel_1_0_15 = pixelVec_1_0_15;
  assign bridge_payload_frame_line_pixel_1_1_0 = pixelVec_1_1_0;
  assign bridge_payload_frame_line_pixel_1_1_1 = pixelVec_1_1_1;
  assign bridge_payload_frame_line_pixel_1_1_2 = pixelVec_1_1_2;
  assign bridge_payload_frame_line_pixel_1_1_3 = pixelVec_1_1_3;
  assign bridge_payload_frame_line_pixel_1_1_4 = pixelVec_1_1_4;
  assign bridge_payload_frame_line_pixel_1_1_5 = pixelVec_1_1_5;
  assign bridge_payload_frame_line_pixel_1_1_6 = pixelVec_1_1_6;
  assign bridge_payload_frame_line_pixel_1_1_7 = pixelVec_1_1_7;
  assign bridge_payload_frame_line_pixel_1_1_8 = pixelVec_1_1_8;
  assign bridge_payload_frame_line_pixel_1_1_9 = pixelVec_1_1_9;
  assign bridge_payload_frame_line_pixel_1_1_10 = pixelVec_1_1_10;
  assign bridge_payload_frame_line_pixel_1_1_11 = pixelVec_1_1_11;
  assign bridge_payload_frame_line_pixel_1_1_12 = pixelVec_1_1_12;
  assign bridge_payload_frame_line_pixel_1_1_13 = pixelVec_1_1_13;
  assign bridge_payload_frame_line_pixel_1_1_14 = pixelVec_1_1_14;
  assign bridge_payload_frame_line_pixel_1_1_15 = pixelVec_1_1_15;
  assign bridge_payload_frame_line_pixel_1_2_0 = pixelVec_1_2_0;
  assign bridge_payload_frame_line_pixel_1_2_1 = pixelVec_1_2_1;
  assign bridge_payload_frame_line_pixel_1_2_2 = pixelVec_1_2_2;
  assign bridge_payload_frame_line_pixel_1_2_3 = pixelVec_1_2_3;
  assign bridge_payload_frame_line_pixel_1_2_4 = pixelVec_1_2_4;
  assign bridge_payload_frame_line_pixel_1_2_5 = pixelVec_1_2_5;
  assign bridge_payload_frame_line_pixel_1_2_6 = pixelVec_1_2_6;
  assign bridge_payload_frame_line_pixel_1_2_7 = pixelVec_1_2_7;
  assign bridge_payload_frame_line_pixel_1_2_8 = pixelVec_1_2_8;
  assign bridge_payload_frame_line_pixel_1_2_9 = pixelVec_1_2_9;
  assign bridge_payload_frame_line_pixel_1_2_10 = pixelVec_1_2_10;
  assign bridge_payload_frame_line_pixel_1_2_11 = pixelVec_1_2_11;
  assign bridge_payload_frame_line_pixel_1_2_12 = pixelVec_1_2_12;
  assign bridge_payload_frame_line_pixel_1_2_13 = pixelVec_1_2_13;
  assign bridge_payload_frame_line_pixel_1_2_14 = pixelVec_1_2_14;
  assign bridge_payload_frame_line_pixel_1_2_15 = pixelVec_1_2_15;
  assign bridge_payload_frame_line_pixel_2_0_0 = down_0_0_0;
  assign bridge_payload_frame_line_pixel_2_0_1 = down_0_0_1;
  assign bridge_payload_frame_line_pixel_2_0_2 = down_0_0_2;
  assign bridge_payload_frame_line_pixel_2_0_3 = down_0_0_3;
  assign bridge_payload_frame_line_pixel_2_0_4 = down_0_0_4;
  assign bridge_payload_frame_line_pixel_2_0_5 = down_0_0_5;
  assign bridge_payload_frame_line_pixel_2_0_6 = down_0_0_6;
  assign bridge_payload_frame_line_pixel_2_0_7 = down_0_0_7;
  assign bridge_payload_frame_line_pixel_2_0_8 = down_0_0_8;
  assign bridge_payload_frame_line_pixel_2_0_9 = down_0_0_9;
  assign bridge_payload_frame_line_pixel_2_0_10 = down_0_0_10;
  assign bridge_payload_frame_line_pixel_2_0_11 = down_0_0_11;
  assign bridge_payload_frame_line_pixel_2_0_12 = down_0_0_12;
  assign bridge_payload_frame_line_pixel_2_0_13 = down_0_0_13;
  assign bridge_payload_frame_line_pixel_2_0_14 = down_0_0_14;
  assign bridge_payload_frame_line_pixel_2_0_15 = down_0_0_15;
  assign bridge_payload_frame_line_pixel_2_1_0 = down_0_1_0;
  assign bridge_payload_frame_line_pixel_2_1_1 = down_0_1_1;
  assign bridge_payload_frame_line_pixel_2_1_2 = down_0_1_2;
  assign bridge_payload_frame_line_pixel_2_1_3 = down_0_1_3;
  assign bridge_payload_frame_line_pixel_2_1_4 = down_0_1_4;
  assign bridge_payload_frame_line_pixel_2_1_5 = down_0_1_5;
  assign bridge_payload_frame_line_pixel_2_1_6 = down_0_1_6;
  assign bridge_payload_frame_line_pixel_2_1_7 = down_0_1_7;
  assign bridge_payload_frame_line_pixel_2_1_8 = down_0_1_8;
  assign bridge_payload_frame_line_pixel_2_1_9 = down_0_1_9;
  assign bridge_payload_frame_line_pixel_2_1_10 = down_0_1_10;
  assign bridge_payload_frame_line_pixel_2_1_11 = down_0_1_11;
  assign bridge_payload_frame_line_pixel_2_1_12 = down_0_1_12;
  assign bridge_payload_frame_line_pixel_2_1_13 = down_0_1_13;
  assign bridge_payload_frame_line_pixel_2_1_14 = down_0_1_14;
  assign bridge_payload_frame_line_pixel_2_1_15 = down_0_1_15;
  assign bridge_payload_frame_line_pixel_2_2_0 = down_0_2_0;
  assign bridge_payload_frame_line_pixel_2_2_1 = down_0_2_1;
  assign bridge_payload_frame_line_pixel_2_2_2 = down_0_2_2;
  assign bridge_payload_frame_line_pixel_2_2_3 = down_0_2_3;
  assign bridge_payload_frame_line_pixel_2_2_4 = down_0_2_4;
  assign bridge_payload_frame_line_pixel_2_2_5 = down_0_2_5;
  assign bridge_payload_frame_line_pixel_2_2_6 = down_0_2_6;
  assign bridge_payload_frame_line_pixel_2_2_7 = down_0_2_7;
  assign bridge_payload_frame_line_pixel_2_2_8 = down_0_2_8;
  assign bridge_payload_frame_line_pixel_2_2_9 = down_0_2_9;
  assign bridge_payload_frame_line_pixel_2_2_10 = down_0_2_10;
  assign bridge_payload_frame_line_pixel_2_2_11 = down_0_2_11;
  assign bridge_payload_frame_line_pixel_2_2_12 = down_0_2_12;
  assign bridge_payload_frame_line_pixel_2_2_13 = down_0_2_13;
  assign bridge_payload_frame_line_pixel_2_2_14 = down_0_2_14;
  assign bridge_payload_frame_line_pixel_2_2_15 = down_0_2_15;
  always @(*) begin
    cnt_willIncrement = 1'b0;
    if(when_PixelBufferSame_l93) begin
      cnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    cnt_willClear = 1'b0;
    if(when_PixelBufferSame_l92) begin
      cnt_willClear = 1'b1;
    end
  end

  assign cnt_willOverflowIfInc = (cnt_value == 1'b1);
  assign cnt_willOverflow = (cnt_willOverflowIfInc && cnt_willIncrement);
  always @(*) begin
    cnt_valueNext = (cnt_value + cnt_willIncrement);
    if(cnt_willClear) begin
      cnt_valueNext = 1'b0;
    end
  end

  assign cntWontOverflowIfInc = (! cnt_willOverflowIfInc);
  assign when_PixelBufferSame_l92 = (bridgeFire && bridge_payload_endOfPack);
  assign when_PixelBufferSame_l93 = (bridgeFire && cntWontOverflowIfInc);
  always @(*) begin
    tmp_videoOut_valid = bridge_valid;
    if(cntWontOverflowIfInc) begin
      tmp_videoOut_valid = 1'b0;
    end
  end

  always @(*) begin
    bridge_ready = videoOut_ready;
    if(cntWontOverflowIfInc) begin
      bridge_ready = 1'b1;
    end
  end

  assign videoOut_valid = tmp_videoOut_valid;
  assign videoOut_payload_frame_line_pixel_0_0_0 = bridge_payload_frame_line_pixel_0_0_0;
  assign videoOut_payload_frame_line_pixel_0_0_1 = bridge_payload_frame_line_pixel_0_0_1;
  assign videoOut_payload_frame_line_pixel_0_0_2 = bridge_payload_frame_line_pixel_0_0_2;
  assign videoOut_payload_frame_line_pixel_0_0_3 = bridge_payload_frame_line_pixel_0_0_3;
  assign videoOut_payload_frame_line_pixel_0_0_4 = bridge_payload_frame_line_pixel_0_0_4;
  assign videoOut_payload_frame_line_pixel_0_0_5 = bridge_payload_frame_line_pixel_0_0_5;
  assign videoOut_payload_frame_line_pixel_0_0_6 = bridge_payload_frame_line_pixel_0_0_6;
  assign videoOut_payload_frame_line_pixel_0_0_7 = bridge_payload_frame_line_pixel_0_0_7;
  assign videoOut_payload_frame_line_pixel_0_0_8 = bridge_payload_frame_line_pixel_0_0_8;
  assign videoOut_payload_frame_line_pixel_0_0_9 = bridge_payload_frame_line_pixel_0_0_9;
  assign videoOut_payload_frame_line_pixel_0_0_10 = bridge_payload_frame_line_pixel_0_0_10;
  assign videoOut_payload_frame_line_pixel_0_0_11 = bridge_payload_frame_line_pixel_0_0_11;
  assign videoOut_payload_frame_line_pixel_0_0_12 = bridge_payload_frame_line_pixel_0_0_12;
  assign videoOut_payload_frame_line_pixel_0_0_13 = bridge_payload_frame_line_pixel_0_0_13;
  assign videoOut_payload_frame_line_pixel_0_0_14 = bridge_payload_frame_line_pixel_0_0_14;
  assign videoOut_payload_frame_line_pixel_0_0_15 = bridge_payload_frame_line_pixel_0_0_15;
  assign videoOut_payload_frame_line_pixel_0_1_0 = bridge_payload_frame_line_pixel_0_1_0;
  assign videoOut_payload_frame_line_pixel_0_1_1 = bridge_payload_frame_line_pixel_0_1_1;
  assign videoOut_payload_frame_line_pixel_0_1_2 = bridge_payload_frame_line_pixel_0_1_2;
  assign videoOut_payload_frame_line_pixel_0_1_3 = bridge_payload_frame_line_pixel_0_1_3;
  assign videoOut_payload_frame_line_pixel_0_1_4 = bridge_payload_frame_line_pixel_0_1_4;
  assign videoOut_payload_frame_line_pixel_0_1_5 = bridge_payload_frame_line_pixel_0_1_5;
  assign videoOut_payload_frame_line_pixel_0_1_6 = bridge_payload_frame_line_pixel_0_1_6;
  assign videoOut_payload_frame_line_pixel_0_1_7 = bridge_payload_frame_line_pixel_0_1_7;
  assign videoOut_payload_frame_line_pixel_0_1_8 = bridge_payload_frame_line_pixel_0_1_8;
  assign videoOut_payload_frame_line_pixel_0_1_9 = bridge_payload_frame_line_pixel_0_1_9;
  assign videoOut_payload_frame_line_pixel_0_1_10 = bridge_payload_frame_line_pixel_0_1_10;
  assign videoOut_payload_frame_line_pixel_0_1_11 = bridge_payload_frame_line_pixel_0_1_11;
  assign videoOut_payload_frame_line_pixel_0_1_12 = bridge_payload_frame_line_pixel_0_1_12;
  assign videoOut_payload_frame_line_pixel_0_1_13 = bridge_payload_frame_line_pixel_0_1_13;
  assign videoOut_payload_frame_line_pixel_0_1_14 = bridge_payload_frame_line_pixel_0_1_14;
  assign videoOut_payload_frame_line_pixel_0_1_15 = bridge_payload_frame_line_pixel_0_1_15;
  assign videoOut_payload_frame_line_pixel_0_2_0 = bridge_payload_frame_line_pixel_0_2_0;
  assign videoOut_payload_frame_line_pixel_0_2_1 = bridge_payload_frame_line_pixel_0_2_1;
  assign videoOut_payload_frame_line_pixel_0_2_2 = bridge_payload_frame_line_pixel_0_2_2;
  assign videoOut_payload_frame_line_pixel_0_2_3 = bridge_payload_frame_line_pixel_0_2_3;
  assign videoOut_payload_frame_line_pixel_0_2_4 = bridge_payload_frame_line_pixel_0_2_4;
  assign videoOut_payload_frame_line_pixel_0_2_5 = bridge_payload_frame_line_pixel_0_2_5;
  assign videoOut_payload_frame_line_pixel_0_2_6 = bridge_payload_frame_line_pixel_0_2_6;
  assign videoOut_payload_frame_line_pixel_0_2_7 = bridge_payload_frame_line_pixel_0_2_7;
  assign videoOut_payload_frame_line_pixel_0_2_8 = bridge_payload_frame_line_pixel_0_2_8;
  assign videoOut_payload_frame_line_pixel_0_2_9 = bridge_payload_frame_line_pixel_0_2_9;
  assign videoOut_payload_frame_line_pixel_0_2_10 = bridge_payload_frame_line_pixel_0_2_10;
  assign videoOut_payload_frame_line_pixel_0_2_11 = bridge_payload_frame_line_pixel_0_2_11;
  assign videoOut_payload_frame_line_pixel_0_2_12 = bridge_payload_frame_line_pixel_0_2_12;
  assign videoOut_payload_frame_line_pixel_0_2_13 = bridge_payload_frame_line_pixel_0_2_13;
  assign videoOut_payload_frame_line_pixel_0_2_14 = bridge_payload_frame_line_pixel_0_2_14;
  assign videoOut_payload_frame_line_pixel_0_2_15 = bridge_payload_frame_line_pixel_0_2_15;
  assign videoOut_payload_frame_line_pixel_1_0_0 = bridge_payload_frame_line_pixel_1_0_0;
  assign videoOut_payload_frame_line_pixel_1_0_1 = bridge_payload_frame_line_pixel_1_0_1;
  assign videoOut_payload_frame_line_pixel_1_0_2 = bridge_payload_frame_line_pixel_1_0_2;
  assign videoOut_payload_frame_line_pixel_1_0_3 = bridge_payload_frame_line_pixel_1_0_3;
  assign videoOut_payload_frame_line_pixel_1_0_4 = bridge_payload_frame_line_pixel_1_0_4;
  assign videoOut_payload_frame_line_pixel_1_0_5 = bridge_payload_frame_line_pixel_1_0_5;
  assign videoOut_payload_frame_line_pixel_1_0_6 = bridge_payload_frame_line_pixel_1_0_6;
  assign videoOut_payload_frame_line_pixel_1_0_7 = bridge_payload_frame_line_pixel_1_0_7;
  assign videoOut_payload_frame_line_pixel_1_0_8 = bridge_payload_frame_line_pixel_1_0_8;
  assign videoOut_payload_frame_line_pixel_1_0_9 = bridge_payload_frame_line_pixel_1_0_9;
  assign videoOut_payload_frame_line_pixel_1_0_10 = bridge_payload_frame_line_pixel_1_0_10;
  assign videoOut_payload_frame_line_pixel_1_0_11 = bridge_payload_frame_line_pixel_1_0_11;
  assign videoOut_payload_frame_line_pixel_1_0_12 = bridge_payload_frame_line_pixel_1_0_12;
  assign videoOut_payload_frame_line_pixel_1_0_13 = bridge_payload_frame_line_pixel_1_0_13;
  assign videoOut_payload_frame_line_pixel_1_0_14 = bridge_payload_frame_line_pixel_1_0_14;
  assign videoOut_payload_frame_line_pixel_1_0_15 = bridge_payload_frame_line_pixel_1_0_15;
  assign videoOut_payload_frame_line_pixel_1_1_0 = bridge_payload_frame_line_pixel_1_1_0;
  assign videoOut_payload_frame_line_pixel_1_1_1 = bridge_payload_frame_line_pixel_1_1_1;
  assign videoOut_payload_frame_line_pixel_1_1_2 = bridge_payload_frame_line_pixel_1_1_2;
  assign videoOut_payload_frame_line_pixel_1_1_3 = bridge_payload_frame_line_pixel_1_1_3;
  assign videoOut_payload_frame_line_pixel_1_1_4 = bridge_payload_frame_line_pixel_1_1_4;
  assign videoOut_payload_frame_line_pixel_1_1_5 = bridge_payload_frame_line_pixel_1_1_5;
  assign videoOut_payload_frame_line_pixel_1_1_6 = bridge_payload_frame_line_pixel_1_1_6;
  assign videoOut_payload_frame_line_pixel_1_1_7 = bridge_payload_frame_line_pixel_1_1_7;
  assign videoOut_payload_frame_line_pixel_1_1_8 = bridge_payload_frame_line_pixel_1_1_8;
  assign videoOut_payload_frame_line_pixel_1_1_9 = bridge_payload_frame_line_pixel_1_1_9;
  assign videoOut_payload_frame_line_pixel_1_1_10 = bridge_payload_frame_line_pixel_1_1_10;
  assign videoOut_payload_frame_line_pixel_1_1_11 = bridge_payload_frame_line_pixel_1_1_11;
  assign videoOut_payload_frame_line_pixel_1_1_12 = bridge_payload_frame_line_pixel_1_1_12;
  assign videoOut_payload_frame_line_pixel_1_1_13 = bridge_payload_frame_line_pixel_1_1_13;
  assign videoOut_payload_frame_line_pixel_1_1_14 = bridge_payload_frame_line_pixel_1_1_14;
  assign videoOut_payload_frame_line_pixel_1_1_15 = bridge_payload_frame_line_pixel_1_1_15;
  assign videoOut_payload_frame_line_pixel_1_2_0 = bridge_payload_frame_line_pixel_1_2_0;
  assign videoOut_payload_frame_line_pixel_1_2_1 = bridge_payload_frame_line_pixel_1_2_1;
  assign videoOut_payload_frame_line_pixel_1_2_2 = bridge_payload_frame_line_pixel_1_2_2;
  assign videoOut_payload_frame_line_pixel_1_2_3 = bridge_payload_frame_line_pixel_1_2_3;
  assign videoOut_payload_frame_line_pixel_1_2_4 = bridge_payload_frame_line_pixel_1_2_4;
  assign videoOut_payload_frame_line_pixel_1_2_5 = bridge_payload_frame_line_pixel_1_2_5;
  assign videoOut_payload_frame_line_pixel_1_2_6 = bridge_payload_frame_line_pixel_1_2_6;
  assign videoOut_payload_frame_line_pixel_1_2_7 = bridge_payload_frame_line_pixel_1_2_7;
  assign videoOut_payload_frame_line_pixel_1_2_8 = bridge_payload_frame_line_pixel_1_2_8;
  assign videoOut_payload_frame_line_pixel_1_2_9 = bridge_payload_frame_line_pixel_1_2_9;
  assign videoOut_payload_frame_line_pixel_1_2_10 = bridge_payload_frame_line_pixel_1_2_10;
  assign videoOut_payload_frame_line_pixel_1_2_11 = bridge_payload_frame_line_pixel_1_2_11;
  assign videoOut_payload_frame_line_pixel_1_2_12 = bridge_payload_frame_line_pixel_1_2_12;
  assign videoOut_payload_frame_line_pixel_1_2_13 = bridge_payload_frame_line_pixel_1_2_13;
  assign videoOut_payload_frame_line_pixel_1_2_14 = bridge_payload_frame_line_pixel_1_2_14;
  assign videoOut_payload_frame_line_pixel_1_2_15 = bridge_payload_frame_line_pixel_1_2_15;
  assign videoOut_payload_frame_line_pixel_2_0_0 = bridge_payload_frame_line_pixel_2_0_0;
  assign videoOut_payload_frame_line_pixel_2_0_1 = bridge_payload_frame_line_pixel_2_0_1;
  assign videoOut_payload_frame_line_pixel_2_0_2 = bridge_payload_frame_line_pixel_2_0_2;
  assign videoOut_payload_frame_line_pixel_2_0_3 = bridge_payload_frame_line_pixel_2_0_3;
  assign videoOut_payload_frame_line_pixel_2_0_4 = bridge_payload_frame_line_pixel_2_0_4;
  assign videoOut_payload_frame_line_pixel_2_0_5 = bridge_payload_frame_line_pixel_2_0_5;
  assign videoOut_payload_frame_line_pixel_2_0_6 = bridge_payload_frame_line_pixel_2_0_6;
  assign videoOut_payload_frame_line_pixel_2_0_7 = bridge_payload_frame_line_pixel_2_0_7;
  assign videoOut_payload_frame_line_pixel_2_0_8 = bridge_payload_frame_line_pixel_2_0_8;
  assign videoOut_payload_frame_line_pixel_2_0_9 = bridge_payload_frame_line_pixel_2_0_9;
  assign videoOut_payload_frame_line_pixel_2_0_10 = bridge_payload_frame_line_pixel_2_0_10;
  assign videoOut_payload_frame_line_pixel_2_0_11 = bridge_payload_frame_line_pixel_2_0_11;
  assign videoOut_payload_frame_line_pixel_2_0_12 = bridge_payload_frame_line_pixel_2_0_12;
  assign videoOut_payload_frame_line_pixel_2_0_13 = bridge_payload_frame_line_pixel_2_0_13;
  assign videoOut_payload_frame_line_pixel_2_0_14 = bridge_payload_frame_line_pixel_2_0_14;
  assign videoOut_payload_frame_line_pixel_2_0_15 = bridge_payload_frame_line_pixel_2_0_15;
  assign videoOut_payload_frame_line_pixel_2_1_0 = bridge_payload_frame_line_pixel_2_1_0;
  assign videoOut_payload_frame_line_pixel_2_1_1 = bridge_payload_frame_line_pixel_2_1_1;
  assign videoOut_payload_frame_line_pixel_2_1_2 = bridge_payload_frame_line_pixel_2_1_2;
  assign videoOut_payload_frame_line_pixel_2_1_3 = bridge_payload_frame_line_pixel_2_1_3;
  assign videoOut_payload_frame_line_pixel_2_1_4 = bridge_payload_frame_line_pixel_2_1_4;
  assign videoOut_payload_frame_line_pixel_2_1_5 = bridge_payload_frame_line_pixel_2_1_5;
  assign videoOut_payload_frame_line_pixel_2_1_6 = bridge_payload_frame_line_pixel_2_1_6;
  assign videoOut_payload_frame_line_pixel_2_1_7 = bridge_payload_frame_line_pixel_2_1_7;
  assign videoOut_payload_frame_line_pixel_2_1_8 = bridge_payload_frame_line_pixel_2_1_8;
  assign videoOut_payload_frame_line_pixel_2_1_9 = bridge_payload_frame_line_pixel_2_1_9;
  assign videoOut_payload_frame_line_pixel_2_1_10 = bridge_payload_frame_line_pixel_2_1_10;
  assign videoOut_payload_frame_line_pixel_2_1_11 = bridge_payload_frame_line_pixel_2_1_11;
  assign videoOut_payload_frame_line_pixel_2_1_12 = bridge_payload_frame_line_pixel_2_1_12;
  assign videoOut_payload_frame_line_pixel_2_1_13 = bridge_payload_frame_line_pixel_2_1_13;
  assign videoOut_payload_frame_line_pixel_2_1_14 = bridge_payload_frame_line_pixel_2_1_14;
  assign videoOut_payload_frame_line_pixel_2_1_15 = bridge_payload_frame_line_pixel_2_1_15;
  assign videoOut_payload_frame_line_pixel_2_2_0 = bridge_payload_frame_line_pixel_2_2_0;
  assign videoOut_payload_frame_line_pixel_2_2_1 = bridge_payload_frame_line_pixel_2_2_1;
  assign videoOut_payload_frame_line_pixel_2_2_2 = bridge_payload_frame_line_pixel_2_2_2;
  assign videoOut_payload_frame_line_pixel_2_2_3 = bridge_payload_frame_line_pixel_2_2_3;
  assign videoOut_payload_frame_line_pixel_2_2_4 = bridge_payload_frame_line_pixel_2_2_4;
  assign videoOut_payload_frame_line_pixel_2_2_5 = bridge_payload_frame_line_pixel_2_2_5;
  assign videoOut_payload_frame_line_pixel_2_2_6 = bridge_payload_frame_line_pixel_2_2_6;
  assign videoOut_payload_frame_line_pixel_2_2_7 = bridge_payload_frame_line_pixel_2_2_7;
  assign videoOut_payload_frame_line_pixel_2_2_8 = bridge_payload_frame_line_pixel_2_2_8;
  assign videoOut_payload_frame_line_pixel_2_2_9 = bridge_payload_frame_line_pixel_2_2_9;
  assign videoOut_payload_frame_line_pixel_2_2_10 = bridge_payload_frame_line_pixel_2_2_10;
  assign videoOut_payload_frame_line_pixel_2_2_11 = bridge_payload_frame_line_pixel_2_2_11;
  assign videoOut_payload_frame_line_pixel_2_2_12 = bridge_payload_frame_line_pixel_2_2_12;
  assign videoOut_payload_frame_line_pixel_2_2_13 = bridge_payload_frame_line_pixel_2_2_13;
  assign videoOut_payload_frame_line_pixel_2_2_14 = bridge_payload_frame_line_pixel_2_2_14;
  assign videoOut_payload_frame_line_pixel_2_2_15 = bridge_payload_frame_line_pixel_2_2_15;
  assign videoOut_payload_frame_line_endOfLine = bridge_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_endOfFrame = bridge_payload_frame_endOfFrame;
  assign videoOut_payload_endOfPack = bridge_payload_endOfPack;
  always @(posedge clk) begin
    if(reset) begin
      paddedCond <= 1'b0;
      cntPrev <= 2'b01;
      cntPost <= 2'b00;
      padded_payload_frame_endOfFrame_delay_1 <= 1'b0;
      padded_payload_frame_line_endOfLine_delay_1 <= 1'b0;
      cnt_value <= 1'b0;
    end else begin
      if(when_PixelBufferSame_l46) begin
        paddedCond <= 1'b1;
      end
      if(tmp_bridge_payload_endOfPack_2) begin
        paddedCond <= 1'b0;
      end
      if(when_PixelBufferSame_l74) begin
        cntPrev <= 2'b00;
      end
      if(when_PixelBufferSame_l75) begin
        cntPost <= 2'b00;
      end
      if(when_PixelBufferSame_l76) begin
        cntPrev <= (cntPrev + 2'b01);
      end
      if(when_PixelBufferSame_l77) begin
        cntPost <= (cntPost + 2'b01);
      end
      if(paddedFire) begin
        padded_payload_frame_endOfFrame_delay_1 <= padded_payload_frame_endOfFrame;
      end
      if(paddedFire) begin
        padded_payload_frame_line_endOfLine_delay_1 <= padded_payload_frame_line_endOfLine;
      end
      cnt_value <= cnt_valueNext;
    end
  end

  always @(posedge clk) begin
    if(paddedFire) begin
      pixelBuffer <= {{{padded_payload_frame_line_pixel_2_15,{padded_payload_frame_line_pixel_2_14,{padded_payload_frame_line_pixel_2_13,{padded_payload_frame_line_pixel_2_12,{tmp_pixelBuffer,tmp_pixelBuffer_1}}}}},{{padded_payload_frame_line_pixel_1_15,{padded_payload_frame_line_pixel_1_14,{padded_payload_frame_line_pixel_1_13,{tmp_pixelBuffer_4,tmp_pixelBuffer_5}}}},{padded_payload_frame_line_pixel_0_15,{padded_payload_frame_line_pixel_0_14,{padded_payload_frame_line_pixel_0_13,{tmp_pixelBuffer_8,tmp_pixelBuffer_9}}}}}},tmp_pixelBuffer_12};
    end
  end


endmodule

module LineBufferSame (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_2_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 videoIn_fork_io_outputs_0_ready;
  reg                 videoIn_fork_io_outputs_1_ready;
  reg                 fifo_pop_fork_io_outputs_0_ready;
  reg                 fifo_pop_fork_io_outputs_1_ready;
  wire                fifo_push_ready;
  wire                fifo_pop_valid;
  wire       [7:0]    fifo_pop_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_payload_0_pixel_15;
  wire                fifo_pop_payload_0_endOfLine;
  wire       [7:0]    fifo_pop_payload_1_pixel_0;
  wire       [7:0]    fifo_pop_payload_1_pixel_1;
  wire       [7:0]    fifo_pop_payload_1_pixel_2;
  wire       [7:0]    fifo_pop_payload_1_pixel_3;
  wire       [7:0]    fifo_pop_payload_1_pixel_4;
  wire       [7:0]    fifo_pop_payload_1_pixel_5;
  wire       [7:0]    fifo_pop_payload_1_pixel_6;
  wire       [7:0]    fifo_pop_payload_1_pixel_7;
  wire       [7:0]    fifo_pop_payload_1_pixel_8;
  wire       [7:0]    fifo_pop_payload_1_pixel_9;
  wire       [7:0]    fifo_pop_payload_1_pixel_10;
  wire       [7:0]    fifo_pop_payload_1_pixel_11;
  wire       [7:0]    fifo_pop_payload_1_pixel_12;
  wire       [7:0]    fifo_pop_payload_1_pixel_13;
  wire       [7:0]    fifo_pop_payload_1_pixel_14;
  wire       [7:0]    fifo_pop_payload_1_pixel_15;
  wire                fifo_pop_payload_1_endOfLine;
  wire                videoIn_fork_io_input_ready;
  wire                videoIn_fork_io_outputs_0_valid;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_0;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_1;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_2;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_3;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_4;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_5;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_6;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_7;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_8;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_9;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_10;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_11;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_12;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_13;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_14;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_15;
  wire                videoIn_fork_io_outputs_0_payload_frame_line_endOfLine;
  wire                videoIn_fork_io_outputs_0_payload_frame_endOfFrame;
  wire                videoIn_fork_io_outputs_0_payload_endOfPack;
  wire                videoIn_fork_io_outputs_1_valid;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_0;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_1;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_2;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_3;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_4;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_5;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_6;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_7;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_8;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_9;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_10;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_11;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_12;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_13;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_14;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_15;
  wire                videoIn_fork_io_outputs_1_payload_frame_line_endOfLine;
  wire                videoIn_fork_io_outputs_1_payload_frame_endOfFrame;
  wire                videoIn_fork_io_outputs_1_payload_endOfPack;
  wire                fifo_pop_fork_io_input_ready;
  wire                fifo_pop_fork_io_outputs_0_valid;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_15;
  wire                fifo_pop_fork_io_outputs_0_payload_0_endOfLine;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_1_pixel_15;
  wire                fifo_pop_fork_io_outputs_0_payload_1_endOfLine;
  wire                fifo_pop_fork_io_outputs_1_valid;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_15;
  wire                fifo_pop_fork_io_outputs_1_payload_0_endOfLine;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_1_pixel_15;
  wire                fifo_pop_fork_io_outputs_1_payload_1_endOfLine;
  wire       [7:0]    zero_0;
  wire       [7:0]    zero_1;
  wire       [7:0]    zero_2;
  wire       [7:0]    zero_3;
  wire       [7:0]    zero_4;
  wire       [7:0]    zero_5;
  wire       [7:0]    zero_6;
  wire       [7:0]    zero_7;
  wire       [7:0]    zero_8;
  wire       [7:0]    zero_9;
  wire       [7:0]    zero_10;
  wire       [7:0]    zero_11;
  wire       [7:0]    zero_12;
  wire       [7:0]    zero_13;
  wire       [7:0]    zero_14;
  wire       [7:0]    zero_15;
  wire       [127:0]  tmp_zero_0;
  wire                in2outThrowCond;
  wire                in2outAddCond;
  wire                in2fifoAddCond;
  wire                fifo2outThrowCond;
  wire                feedbackThrowCond;
  wire                feedbackAddCond;
  reg                 tmp_in2outThrownAdded_valid;
  reg                 tmp_io_outputs_1_ready;
  reg                 in2outThrownAdded_valid;
  wire                in2outThrownAdded_ready;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_0;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_1;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_2;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_3;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_4;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_5;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_6;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_7;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_8;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_9;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_10;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_11;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_12;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_13;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_14;
  wire       [7:0]    in2outThrownAdded_payload_frame_line_pixel_15;
  wire                in2outThrownAdded_payload_frame_line_endOfLine;
  wire                in2outThrownAdded_payload_frame_endOfFrame;
  wire                in2outThrownAdded_payload_endOfPack;
  reg                 in2fifoAdded_valid;
  wire                in2fifoAdded_ready;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_0;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_1;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_2;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_3;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_4;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_5;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_6;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_7;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_8;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_9;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_10;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_11;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_12;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_13;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_14;
  wire       [7:0]    in2fifoAdded_payload_frame_line_pixel_15;
  wire                in2fifoAdded_payload_frame_line_endOfLine;
  wire                in2fifoAdded_payload_frame_endOfFrame;
  wire                in2fifoAdded_payload_endOfPack;
  reg                 fifo2outThrown_valid;
  wire                fifo2outThrown_ready;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_0;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_1;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_2;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_3;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_4;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_5;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_6;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_7;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_8;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_9;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_10;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_11;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_12;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_13;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_14;
  wire       [7:0]    fifo2outThrown_payload_0_pixel_15;
  wire                fifo2outThrown_payload_0_endOfLine;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_0;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_1;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_2;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_3;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_4;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_5;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_6;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_7;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_8;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_9;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_10;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_11;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_12;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_13;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_14;
  wire       [7:0]    fifo2outThrown_payload_1_pixel_15;
  wire                fifo2outThrown_payload_1_endOfLine;
  reg                 tmp_feedbackThrownAdded_valid;
  reg                 tmp_io_outputs_0_ready;
  reg                 feedbackThrownAdded_valid;
  wire                feedbackThrownAdded_ready;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_0;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_1;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_2;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_3;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_4;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_5;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_6;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_7;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_8;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_9;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_10;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_11;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_12;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_13;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_14;
  wire       [7:0]    feedbackThrownAdded_payload_0_pixel_15;
  wire                feedbackThrownAdded_payload_0_endOfLine;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_0;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_1;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_2;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_3;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_4;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_5;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_6;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_7;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_8;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_9;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_10;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_11;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_12;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_13;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_14;
  wire       [7:0]    feedbackThrownAdded_payload_1_pixel_15;
  wire                feedbackThrownAdded_payload_1_endOfLine;
  wire                in2fifoJoinFeedback_valid;
  wire                in2fifoJoinFeedback_ready;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_0;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_1;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_2;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_3;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_4;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_5;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_6;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_7;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_8;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_9;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_10;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_11;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_12;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_13;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_14;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_15;
  wire                in2fifoJoinFeedback_payload__1_frame_line_endOfLine;
  wire                in2fifoJoinFeedback_payload__1_frame_endOfFrame;
  wire                in2fifoJoinFeedback_payload__1_endOfPack;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_0;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_1;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_2;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_3;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_4;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_5;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_6;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_7;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_8;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_9;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_10;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_11;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_12;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_13;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_14;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_15;
  wire                in2fifoJoinFeedback_payload__2_0_endOfLine;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_0;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_1;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_2;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_3;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_4;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_5;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_6;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_7;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_8;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_9;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_10;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_11;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_12;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_13;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_14;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_1_pixel_15;
  wire                in2fifoJoinFeedback_payload__2_1_endOfLine;
  wire                in2fifoJoinFeedback_fire;
  wire                in2fifoJoinFeedback_fire_1;
  wire                in2outJoinFifo2out_valid;
  wire                in2outJoinFifo2out_ready;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_0;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_1;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_2;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_3;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_4;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_5;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_6;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_7;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_8;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_9;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_10;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_11;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_12;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_13;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_14;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_15;
  wire                in2outJoinFifo2out_payload__1_frame_line_endOfLine;
  wire                in2outJoinFifo2out_payload__1_frame_endOfFrame;
  wire                in2outJoinFifo2out_payload__1_endOfPack;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_0;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_1;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_2;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_3;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_4;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_5;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_6;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_7;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_8;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_9;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_10;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_11;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_12;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_13;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_14;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_15;
  wire                in2outJoinFifo2out_payload__2_0_endOfLine;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_0;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_1;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_2;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_3;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_4;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_5;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_6;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_7;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_8;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_9;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_10;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_11;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_12;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_13;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_14;
  wire       [7:0]    in2outJoinFifo2out_payload__2_1_pixel_15;
  wire                in2outJoinFifo2out_payload__2_1_endOfLine;
  wire                in2outJoinFifo2out_fire;
  wire                in2outJoinFifo2out_fire_1;
  reg                 firstFewLines_willIncrement;
  reg                 firstFewLines_willClear;
  reg        [0:0]    firstFewLines_valueNext;
  reg        [0:0]    firstFewLines_value;
  wire                firstFewLines_willOverflowIfInc;
  wire                firstFewLines_willOverflow;
  wire                ioVideoInFire;
  wire                firstLine;
  wire                firstFewLinesWontOverflowIfInc;
  wire                when_LineBufferSame_l71;
  wire                when_LineBufferSame_l72;
  reg                 lastFewLines_willIncrement;
  reg                 lastFewLines_willClear;
  wire                lastFewLines_willOverflowIfInc;
  wire                lastFewLines_willOverflow;
  wire                ioVideoOutFire;
  wire                lastFewLinesWontOverflowIfInc;
  wire                when_LineBufferSame_l77;
  wire                when_LineBufferSame_l78;
  reg                 endOfFrameGap;
  wire                when_LineBufferSame_l81;
  wire                when_LineBufferSame_l81_1;
  reg                 endOfPackGap;
  wire                when_LineBufferSame_l83;
  wire                when_LineBufferSame_l83_1;
  wire                endOfPackGapInv;
  reg        [1:0]    cntPrev;
  reg        [1:0]    cntPost;
  wire                cntPrevStable;
  wire                cntPostStable;
  wire                cntPrevEqualVec_0;
  wire                cntPostEqualVec_0;
  wire                when_LineBufferSame_l103;
  wire                when_LineBufferSame_l104;
  wire                when_LineBufferSame_l105;
  wire                when_LineBufferSame_l106;
  wire       [7:0]    up_0_0;
  wire       [7:0]    up_0_1;
  wire       [7:0]    up_0_2;
  wire       [7:0]    up_0_3;
  wire       [7:0]    up_0_4;
  wire       [7:0]    up_0_5;
  wire       [7:0]    up_0_6;
  wire       [7:0]    up_0_7;
  wire       [7:0]    up_0_8;
  wire       [7:0]    up_0_9;
  wire       [7:0]    up_0_10;
  wire       [7:0]    up_0_11;
  wire       [7:0]    up_0_12;
  wire       [7:0]    up_0_13;
  wire       [7:0]    up_0_14;
  wire       [7:0]    up_0_15;
  wire       [7:0]    down_0_0;
  wire       [7:0]    down_0_1;
  wire       [7:0]    down_0_2;
  wire       [7:0]    down_0_3;
  wire       [7:0]    down_0_4;
  wire       [7:0]    down_0_5;
  wire       [7:0]    down_0_6;
  wire       [7:0]    down_0_7;
  wire       [7:0]    down_0_8;
  wire       [7:0]    down_0_9;
  wire       [7:0]    down_0_10;
  wire       [7:0]    down_0_11;
  wire       [7:0]    down_0_12;
  wire       [7:0]    down_0_13;
  wire       [7:0]    down_0_14;
  wire       [7:0]    down_0_15;

  StreamFifoHighPerf_1 fifo (
    .push_valid                  (in2fifoJoinFeedback_valid                                ), //i
    .push_ready                  (fifo_push_ready                                          ), //o
    .push_payload_0_pixel_0      (in2fifoJoinFeedback_payload__2_1_pixel_0[7:0]            ), //i
    .push_payload_0_pixel_1      (in2fifoJoinFeedback_payload__2_1_pixel_1[7:0]            ), //i
    .push_payload_0_pixel_2      (in2fifoJoinFeedback_payload__2_1_pixel_2[7:0]            ), //i
    .push_payload_0_pixel_3      (in2fifoJoinFeedback_payload__2_1_pixel_3[7:0]            ), //i
    .push_payload_0_pixel_4      (in2fifoJoinFeedback_payload__2_1_pixel_4[7:0]            ), //i
    .push_payload_0_pixel_5      (in2fifoJoinFeedback_payload__2_1_pixel_5[7:0]            ), //i
    .push_payload_0_pixel_6      (in2fifoJoinFeedback_payload__2_1_pixel_6[7:0]            ), //i
    .push_payload_0_pixel_7      (in2fifoJoinFeedback_payload__2_1_pixel_7[7:0]            ), //i
    .push_payload_0_pixel_8      (in2fifoJoinFeedback_payload__2_1_pixel_8[7:0]            ), //i
    .push_payload_0_pixel_9      (in2fifoJoinFeedback_payload__2_1_pixel_9[7:0]            ), //i
    .push_payload_0_pixel_10     (in2fifoJoinFeedback_payload__2_1_pixel_10[7:0]           ), //i
    .push_payload_0_pixel_11     (in2fifoJoinFeedback_payload__2_1_pixel_11[7:0]           ), //i
    .push_payload_0_pixel_12     (in2fifoJoinFeedback_payload__2_1_pixel_12[7:0]           ), //i
    .push_payload_0_pixel_13     (in2fifoJoinFeedback_payload__2_1_pixel_13[7:0]           ), //i
    .push_payload_0_pixel_14     (in2fifoJoinFeedback_payload__2_1_pixel_14[7:0]           ), //i
    .push_payload_0_pixel_15     (in2fifoJoinFeedback_payload__2_1_pixel_15[7:0]           ), //i
    .push_payload_0_endOfLine    (in2fifoJoinFeedback_payload__2_1_endOfLine               ), //i
    .push_payload_1_pixel_0      (in2fifoJoinFeedback_payload__1_frame_line_pixel_0[7:0]   ), //i
    .push_payload_1_pixel_1      (in2fifoJoinFeedback_payload__1_frame_line_pixel_1[7:0]   ), //i
    .push_payload_1_pixel_2      (in2fifoJoinFeedback_payload__1_frame_line_pixel_2[7:0]   ), //i
    .push_payload_1_pixel_3      (in2fifoJoinFeedback_payload__1_frame_line_pixel_3[7:0]   ), //i
    .push_payload_1_pixel_4      (in2fifoJoinFeedback_payload__1_frame_line_pixel_4[7:0]   ), //i
    .push_payload_1_pixel_5      (in2fifoJoinFeedback_payload__1_frame_line_pixel_5[7:0]   ), //i
    .push_payload_1_pixel_6      (in2fifoJoinFeedback_payload__1_frame_line_pixel_6[7:0]   ), //i
    .push_payload_1_pixel_7      (in2fifoJoinFeedback_payload__1_frame_line_pixel_7[7:0]   ), //i
    .push_payload_1_pixel_8      (in2fifoJoinFeedback_payload__1_frame_line_pixel_8[7:0]   ), //i
    .push_payload_1_pixel_9      (in2fifoJoinFeedback_payload__1_frame_line_pixel_9[7:0]   ), //i
    .push_payload_1_pixel_10     (in2fifoJoinFeedback_payload__1_frame_line_pixel_10[7:0]  ), //i
    .push_payload_1_pixel_11     (in2fifoJoinFeedback_payload__1_frame_line_pixel_11[7:0]  ), //i
    .push_payload_1_pixel_12     (in2fifoJoinFeedback_payload__1_frame_line_pixel_12[7:0]  ), //i
    .push_payload_1_pixel_13     (in2fifoJoinFeedback_payload__1_frame_line_pixel_13[7:0]  ), //i
    .push_payload_1_pixel_14     (in2fifoJoinFeedback_payload__1_frame_line_pixel_14[7:0]  ), //i
    .push_payload_1_pixel_15     (in2fifoJoinFeedback_payload__1_frame_line_pixel_15[7:0]  ), //i
    .push_payload_1_endOfLine    (in2fifoJoinFeedback_payload__1_frame_line_endOfLine      ), //i
    .pop_valid                   (fifo_pop_valid                                           ), //o
    .pop_ready                   (fifo_pop_fork_io_input_ready                             ), //i
    .pop_payload_0_pixel_0       (fifo_pop_payload_0_pixel_0[7:0]                          ), //o
    .pop_payload_0_pixel_1       (fifo_pop_payload_0_pixel_1[7:0]                          ), //o
    .pop_payload_0_pixel_2       (fifo_pop_payload_0_pixel_2[7:0]                          ), //o
    .pop_payload_0_pixel_3       (fifo_pop_payload_0_pixel_3[7:0]                          ), //o
    .pop_payload_0_pixel_4       (fifo_pop_payload_0_pixel_4[7:0]                          ), //o
    .pop_payload_0_pixel_5       (fifo_pop_payload_0_pixel_5[7:0]                          ), //o
    .pop_payload_0_pixel_6       (fifo_pop_payload_0_pixel_6[7:0]                          ), //o
    .pop_payload_0_pixel_7       (fifo_pop_payload_0_pixel_7[7:0]                          ), //o
    .pop_payload_0_pixel_8       (fifo_pop_payload_0_pixel_8[7:0]                          ), //o
    .pop_payload_0_pixel_9       (fifo_pop_payload_0_pixel_9[7:0]                          ), //o
    .pop_payload_0_pixel_10      (fifo_pop_payload_0_pixel_10[7:0]                         ), //o
    .pop_payload_0_pixel_11      (fifo_pop_payload_0_pixel_11[7:0]                         ), //o
    .pop_payload_0_pixel_12      (fifo_pop_payload_0_pixel_12[7:0]                         ), //o
    .pop_payload_0_pixel_13      (fifo_pop_payload_0_pixel_13[7:0]                         ), //o
    .pop_payload_0_pixel_14      (fifo_pop_payload_0_pixel_14[7:0]                         ), //o
    .pop_payload_0_pixel_15      (fifo_pop_payload_0_pixel_15[7:0]                         ), //o
    .pop_payload_0_endOfLine     (fifo_pop_payload_0_endOfLine                             ), //o
    .pop_payload_1_pixel_0       (fifo_pop_payload_1_pixel_0[7:0]                          ), //o
    .pop_payload_1_pixel_1       (fifo_pop_payload_1_pixel_1[7:0]                          ), //o
    .pop_payload_1_pixel_2       (fifo_pop_payload_1_pixel_2[7:0]                          ), //o
    .pop_payload_1_pixel_3       (fifo_pop_payload_1_pixel_3[7:0]                          ), //o
    .pop_payload_1_pixel_4       (fifo_pop_payload_1_pixel_4[7:0]                          ), //o
    .pop_payload_1_pixel_5       (fifo_pop_payload_1_pixel_5[7:0]                          ), //o
    .pop_payload_1_pixel_6       (fifo_pop_payload_1_pixel_6[7:0]                          ), //o
    .pop_payload_1_pixel_7       (fifo_pop_payload_1_pixel_7[7:0]                          ), //o
    .pop_payload_1_pixel_8       (fifo_pop_payload_1_pixel_8[7:0]                          ), //o
    .pop_payload_1_pixel_9       (fifo_pop_payload_1_pixel_9[7:0]                          ), //o
    .pop_payload_1_pixel_10      (fifo_pop_payload_1_pixel_10[7:0]                         ), //o
    .pop_payload_1_pixel_11      (fifo_pop_payload_1_pixel_11[7:0]                         ), //o
    .pop_payload_1_pixel_12      (fifo_pop_payload_1_pixel_12[7:0]                         ), //o
    .pop_payload_1_pixel_13      (fifo_pop_payload_1_pixel_13[7:0]                         ), //o
    .pop_payload_1_pixel_14      (fifo_pop_payload_1_pixel_14[7:0]                         ), //o
    .pop_payload_1_pixel_15      (fifo_pop_payload_1_pixel_15[7:0]                         ), //o
    .pop_payload_1_endOfLine     (fifo_pop_payload_1_endOfLine                             ), //o
    .flush                       (1'b0                                                     ), //i
    .clk                         (clk                                                      ), //i
    .reset                       (reset                                                    )  //i
  );
  StreamFork videoIn_fork (
    .io_input_valid                               (videoIn_valid                                               ), //i
    .io_input_ready                               (videoIn_fork_io_input_ready                                 ), //o
    .io_input_payload_frame_line_pixel_0          (videoIn_payload_frame_line_pixel_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1          (videoIn_payload_frame_line_pixel_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2          (videoIn_payload_frame_line_pixel_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_3          (videoIn_payload_frame_line_pixel_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_4          (videoIn_payload_frame_line_pixel_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_5          (videoIn_payload_frame_line_pixel_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_6          (videoIn_payload_frame_line_pixel_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_7          (videoIn_payload_frame_line_pixel_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_8          (videoIn_payload_frame_line_pixel_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_9          (videoIn_payload_frame_line_pixel_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_10         (videoIn_payload_frame_line_pixel_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_11         (videoIn_payload_frame_line_pixel_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_12         (videoIn_payload_frame_line_pixel_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_13         (videoIn_payload_frame_line_pixel_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_14         (videoIn_payload_frame_line_pixel_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_15         (videoIn_payload_frame_line_pixel_15[7:0]                    ), //i
    .io_input_payload_frame_line_endOfLine        (videoIn_payload_frame_line_endOfLine                        ), //i
    .io_input_payload_frame_endOfFrame            (videoIn_payload_frame_endOfFrame                            ), //i
    .io_input_payload_endOfPack                   (videoIn_payload_endOfPack                                   ), //i
    .io_outputs_0_valid                           (videoIn_fork_io_outputs_0_valid                             ), //o
    .io_outputs_0_ready                           (videoIn_fork_io_outputs_0_ready                             ), //i
    .io_outputs_0_payload_frame_line_pixel_0      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_3      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_4      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_5      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_6      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_7      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_8      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_9      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_10     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_11     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_12     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_13     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_14     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_15     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_endOfLine    (videoIn_fork_io_outputs_0_payload_frame_line_endOfLine      ), //o
    .io_outputs_0_payload_frame_endOfFrame        (videoIn_fork_io_outputs_0_payload_frame_endOfFrame          ), //o
    .io_outputs_0_payload_endOfPack               (videoIn_fork_io_outputs_0_payload_endOfPack                 ), //o
    .io_outputs_1_valid                           (videoIn_fork_io_outputs_1_valid                             ), //o
    .io_outputs_1_ready                           (videoIn_fork_io_outputs_1_ready                             ), //i
    .io_outputs_1_payload_frame_line_pixel_0      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_3      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_4      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_5      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_6      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_7      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_8      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_9      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_10     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_11     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_12     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_13     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_14     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_15     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_endOfLine    (videoIn_fork_io_outputs_1_payload_frame_line_endOfLine      ), //o
    .io_outputs_1_payload_frame_endOfFrame        (videoIn_fork_io_outputs_1_payload_frame_endOfFrame          ), //o
    .io_outputs_1_payload_endOfPack               (videoIn_fork_io_outputs_1_payload_endOfPack                 ), //o
    .clk                                          (clk                                                         ), //i
    .reset                                        (reset                                                       )  //i
  );
  StreamFork_3 fifo_pop_fork (
    .io_input_valid                      (fifo_pop_valid                                      ), //i
    .io_input_ready                      (fifo_pop_fork_io_input_ready                        ), //o
    .io_input_payload_0_pixel_0          (fifo_pop_payload_0_pixel_0[7:0]                     ), //i
    .io_input_payload_0_pixel_1          (fifo_pop_payload_0_pixel_1[7:0]                     ), //i
    .io_input_payload_0_pixel_2          (fifo_pop_payload_0_pixel_2[7:0]                     ), //i
    .io_input_payload_0_pixel_3          (fifo_pop_payload_0_pixel_3[7:0]                     ), //i
    .io_input_payload_0_pixel_4          (fifo_pop_payload_0_pixel_4[7:0]                     ), //i
    .io_input_payload_0_pixel_5          (fifo_pop_payload_0_pixel_5[7:0]                     ), //i
    .io_input_payload_0_pixel_6          (fifo_pop_payload_0_pixel_6[7:0]                     ), //i
    .io_input_payload_0_pixel_7          (fifo_pop_payload_0_pixel_7[7:0]                     ), //i
    .io_input_payload_0_pixel_8          (fifo_pop_payload_0_pixel_8[7:0]                     ), //i
    .io_input_payload_0_pixel_9          (fifo_pop_payload_0_pixel_9[7:0]                     ), //i
    .io_input_payload_0_pixel_10         (fifo_pop_payload_0_pixel_10[7:0]                    ), //i
    .io_input_payload_0_pixel_11         (fifo_pop_payload_0_pixel_11[7:0]                    ), //i
    .io_input_payload_0_pixel_12         (fifo_pop_payload_0_pixel_12[7:0]                    ), //i
    .io_input_payload_0_pixel_13         (fifo_pop_payload_0_pixel_13[7:0]                    ), //i
    .io_input_payload_0_pixel_14         (fifo_pop_payload_0_pixel_14[7:0]                    ), //i
    .io_input_payload_0_pixel_15         (fifo_pop_payload_0_pixel_15[7:0]                    ), //i
    .io_input_payload_0_endOfLine        (fifo_pop_payload_0_endOfLine                        ), //i
    .io_input_payload_1_pixel_0          (fifo_pop_payload_1_pixel_0[7:0]                     ), //i
    .io_input_payload_1_pixel_1          (fifo_pop_payload_1_pixel_1[7:0]                     ), //i
    .io_input_payload_1_pixel_2          (fifo_pop_payload_1_pixel_2[7:0]                     ), //i
    .io_input_payload_1_pixel_3          (fifo_pop_payload_1_pixel_3[7:0]                     ), //i
    .io_input_payload_1_pixel_4          (fifo_pop_payload_1_pixel_4[7:0]                     ), //i
    .io_input_payload_1_pixel_5          (fifo_pop_payload_1_pixel_5[7:0]                     ), //i
    .io_input_payload_1_pixel_6          (fifo_pop_payload_1_pixel_6[7:0]                     ), //i
    .io_input_payload_1_pixel_7          (fifo_pop_payload_1_pixel_7[7:0]                     ), //i
    .io_input_payload_1_pixel_8          (fifo_pop_payload_1_pixel_8[7:0]                     ), //i
    .io_input_payload_1_pixel_9          (fifo_pop_payload_1_pixel_9[7:0]                     ), //i
    .io_input_payload_1_pixel_10         (fifo_pop_payload_1_pixel_10[7:0]                    ), //i
    .io_input_payload_1_pixel_11         (fifo_pop_payload_1_pixel_11[7:0]                    ), //i
    .io_input_payload_1_pixel_12         (fifo_pop_payload_1_pixel_12[7:0]                    ), //i
    .io_input_payload_1_pixel_13         (fifo_pop_payload_1_pixel_13[7:0]                    ), //i
    .io_input_payload_1_pixel_14         (fifo_pop_payload_1_pixel_14[7:0]                    ), //i
    .io_input_payload_1_pixel_15         (fifo_pop_payload_1_pixel_15[7:0]                    ), //i
    .io_input_payload_1_endOfLine        (fifo_pop_payload_1_endOfLine                        ), //i
    .io_outputs_0_valid                  (fifo_pop_fork_io_outputs_0_valid                    ), //o
    .io_outputs_0_ready                  (fifo_pop_fork_io_outputs_0_ready                    ), //i
    .io_outputs_0_payload_0_pixel_0      (fifo_pop_fork_io_outputs_0_payload_0_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_1      (fifo_pop_fork_io_outputs_0_payload_0_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_2      (fifo_pop_fork_io_outputs_0_payload_0_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_3      (fifo_pop_fork_io_outputs_0_payload_0_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_4      (fifo_pop_fork_io_outputs_0_payload_0_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_5      (fifo_pop_fork_io_outputs_0_payload_0_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_6      (fifo_pop_fork_io_outputs_0_payload_0_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_7      (fifo_pop_fork_io_outputs_0_payload_0_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_8      (fifo_pop_fork_io_outputs_0_payload_0_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_9      (fifo_pop_fork_io_outputs_0_payload_0_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_10     (fifo_pop_fork_io_outputs_0_payload_0_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_11     (fifo_pop_fork_io_outputs_0_payload_0_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_12     (fifo_pop_fork_io_outputs_0_payload_0_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_13     (fifo_pop_fork_io_outputs_0_payload_0_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_14     (fifo_pop_fork_io_outputs_0_payload_0_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_15     (fifo_pop_fork_io_outputs_0_payload_0_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_0_endOfLine    (fifo_pop_fork_io_outputs_0_payload_0_endOfLine      ), //o
    .io_outputs_0_payload_1_pixel_0      (fifo_pop_fork_io_outputs_0_payload_1_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_1      (fifo_pop_fork_io_outputs_0_payload_1_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_2      (fifo_pop_fork_io_outputs_0_payload_1_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_3      (fifo_pop_fork_io_outputs_0_payload_1_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_4      (fifo_pop_fork_io_outputs_0_payload_1_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_5      (fifo_pop_fork_io_outputs_0_payload_1_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_6      (fifo_pop_fork_io_outputs_0_payload_1_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_7      (fifo_pop_fork_io_outputs_0_payload_1_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_8      (fifo_pop_fork_io_outputs_0_payload_1_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_9      (fifo_pop_fork_io_outputs_0_payload_1_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_1_pixel_10     (fifo_pop_fork_io_outputs_0_payload_1_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_1_pixel_11     (fifo_pop_fork_io_outputs_0_payload_1_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_1_pixel_12     (fifo_pop_fork_io_outputs_0_payload_1_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_1_pixel_13     (fifo_pop_fork_io_outputs_0_payload_1_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_1_pixel_14     (fifo_pop_fork_io_outputs_0_payload_1_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_1_pixel_15     (fifo_pop_fork_io_outputs_0_payload_1_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_1_endOfLine    (fifo_pop_fork_io_outputs_0_payload_1_endOfLine      ), //o
    .io_outputs_1_valid                  (fifo_pop_fork_io_outputs_1_valid                    ), //o
    .io_outputs_1_ready                  (fifo_pop_fork_io_outputs_1_ready                    ), //i
    .io_outputs_1_payload_0_pixel_0      (fifo_pop_fork_io_outputs_1_payload_0_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_1      (fifo_pop_fork_io_outputs_1_payload_0_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_2      (fifo_pop_fork_io_outputs_1_payload_0_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_3      (fifo_pop_fork_io_outputs_1_payload_0_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_4      (fifo_pop_fork_io_outputs_1_payload_0_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_5      (fifo_pop_fork_io_outputs_1_payload_0_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_6      (fifo_pop_fork_io_outputs_1_payload_0_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_7      (fifo_pop_fork_io_outputs_1_payload_0_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_8      (fifo_pop_fork_io_outputs_1_payload_0_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_9      (fifo_pop_fork_io_outputs_1_payload_0_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_10     (fifo_pop_fork_io_outputs_1_payload_0_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_11     (fifo_pop_fork_io_outputs_1_payload_0_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_12     (fifo_pop_fork_io_outputs_1_payload_0_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_13     (fifo_pop_fork_io_outputs_1_payload_0_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_14     (fifo_pop_fork_io_outputs_1_payload_0_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_15     (fifo_pop_fork_io_outputs_1_payload_0_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_0_endOfLine    (fifo_pop_fork_io_outputs_1_payload_0_endOfLine      ), //o
    .io_outputs_1_payload_1_pixel_0      (fifo_pop_fork_io_outputs_1_payload_1_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_1      (fifo_pop_fork_io_outputs_1_payload_1_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_2      (fifo_pop_fork_io_outputs_1_payload_1_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_3      (fifo_pop_fork_io_outputs_1_payload_1_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_4      (fifo_pop_fork_io_outputs_1_payload_1_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_5      (fifo_pop_fork_io_outputs_1_payload_1_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_6      (fifo_pop_fork_io_outputs_1_payload_1_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_7      (fifo_pop_fork_io_outputs_1_payload_1_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_8      (fifo_pop_fork_io_outputs_1_payload_1_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_9      (fifo_pop_fork_io_outputs_1_payload_1_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_1_pixel_10     (fifo_pop_fork_io_outputs_1_payload_1_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_1_pixel_11     (fifo_pop_fork_io_outputs_1_payload_1_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_1_pixel_12     (fifo_pop_fork_io_outputs_1_payload_1_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_1_pixel_13     (fifo_pop_fork_io_outputs_1_payload_1_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_1_pixel_14     (fifo_pop_fork_io_outputs_1_payload_1_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_1_pixel_15     (fifo_pop_fork_io_outputs_1_payload_1_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_1_endOfLine    (fifo_pop_fork_io_outputs_1_payload_1_endOfLine      ), //o
    .clk                                 (clk                                                 ), //i
    .reset                               (reset                                               )  //i
  );
  assign tmp_zero_0 = 128'h0;
  assign zero_0 = tmp_zero_0[7 : 0];
  assign zero_1 = tmp_zero_0[15 : 8];
  assign zero_2 = tmp_zero_0[23 : 16];
  assign zero_3 = tmp_zero_0[31 : 24];
  assign zero_4 = tmp_zero_0[39 : 32];
  assign zero_5 = tmp_zero_0[47 : 40];
  assign zero_6 = tmp_zero_0[55 : 48];
  assign zero_7 = tmp_zero_0[63 : 56];
  assign zero_8 = tmp_zero_0[71 : 64];
  assign zero_9 = tmp_zero_0[79 : 72];
  assign zero_10 = tmp_zero_0[87 : 80];
  assign zero_11 = tmp_zero_0[95 : 88];
  assign zero_12 = tmp_zero_0[103 : 96];
  assign zero_13 = tmp_zero_0[111 : 104];
  assign zero_14 = tmp_zero_0[119 : 112];
  assign zero_15 = tmp_zero_0[127 : 120];
  assign videoIn_ready = videoIn_fork_io_input_ready;
  always @(*) begin
    tmp_in2outThrownAdded_valid = videoIn_fork_io_outputs_1_valid;
    if(in2outThrowCond) begin
      tmp_in2outThrownAdded_valid = 1'b0;
    end
  end

  always @(*) begin
    videoIn_fork_io_outputs_1_ready = tmp_io_outputs_1_ready;
    if(in2outThrowCond) begin
      videoIn_fork_io_outputs_1_ready = 1'b1;
    end
  end

  always @(*) begin
    in2outThrownAdded_valid = tmp_in2outThrownAdded_valid;
    if(in2outAddCond) begin
      in2outThrownAdded_valid = 1'b1;
    end
  end

  always @(*) begin
    tmp_io_outputs_1_ready = in2outThrownAdded_ready;
    if(in2outAddCond) begin
      tmp_io_outputs_1_ready = 1'b0;
    end
  end

  assign in2outThrownAdded_payload_frame_line_pixel_0 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_0;
  assign in2outThrownAdded_payload_frame_line_pixel_1 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_1;
  assign in2outThrownAdded_payload_frame_line_pixel_2 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_2;
  assign in2outThrownAdded_payload_frame_line_pixel_3 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_3;
  assign in2outThrownAdded_payload_frame_line_pixel_4 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_4;
  assign in2outThrownAdded_payload_frame_line_pixel_5 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_5;
  assign in2outThrownAdded_payload_frame_line_pixel_6 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_6;
  assign in2outThrownAdded_payload_frame_line_pixel_7 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_7;
  assign in2outThrownAdded_payload_frame_line_pixel_8 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_8;
  assign in2outThrownAdded_payload_frame_line_pixel_9 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_9;
  assign in2outThrownAdded_payload_frame_line_pixel_10 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_10;
  assign in2outThrownAdded_payload_frame_line_pixel_11 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_11;
  assign in2outThrownAdded_payload_frame_line_pixel_12 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_12;
  assign in2outThrownAdded_payload_frame_line_pixel_13 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_13;
  assign in2outThrownAdded_payload_frame_line_pixel_14 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_14;
  assign in2outThrownAdded_payload_frame_line_pixel_15 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_15;
  assign in2outThrownAdded_payload_frame_line_endOfLine = videoIn_fork_io_outputs_1_payload_frame_line_endOfLine;
  assign in2outThrownAdded_payload_frame_endOfFrame = videoIn_fork_io_outputs_1_payload_frame_endOfFrame;
  assign in2outThrownAdded_payload_endOfPack = videoIn_fork_io_outputs_1_payload_endOfPack;
  always @(*) begin
    in2fifoAdded_valid = videoIn_fork_io_outputs_0_valid;
    if(in2fifoAddCond) begin
      in2fifoAdded_valid = 1'b1;
    end
  end

  always @(*) begin
    videoIn_fork_io_outputs_0_ready = in2fifoAdded_ready;
    if(in2fifoAddCond) begin
      videoIn_fork_io_outputs_0_ready = 1'b0;
    end
  end

  assign in2fifoAdded_payload_frame_line_pixel_0 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_0;
  assign in2fifoAdded_payload_frame_line_pixel_1 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_1;
  assign in2fifoAdded_payload_frame_line_pixel_2 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_2;
  assign in2fifoAdded_payload_frame_line_pixel_3 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_3;
  assign in2fifoAdded_payload_frame_line_pixel_4 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_4;
  assign in2fifoAdded_payload_frame_line_pixel_5 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_5;
  assign in2fifoAdded_payload_frame_line_pixel_6 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_6;
  assign in2fifoAdded_payload_frame_line_pixel_7 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_7;
  assign in2fifoAdded_payload_frame_line_pixel_8 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_8;
  assign in2fifoAdded_payload_frame_line_pixel_9 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_9;
  assign in2fifoAdded_payload_frame_line_pixel_10 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_10;
  assign in2fifoAdded_payload_frame_line_pixel_11 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_11;
  assign in2fifoAdded_payload_frame_line_pixel_12 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_12;
  assign in2fifoAdded_payload_frame_line_pixel_13 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_13;
  assign in2fifoAdded_payload_frame_line_pixel_14 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_14;
  assign in2fifoAdded_payload_frame_line_pixel_15 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_15;
  assign in2fifoAdded_payload_frame_line_endOfLine = videoIn_fork_io_outputs_0_payload_frame_line_endOfLine;
  assign in2fifoAdded_payload_frame_endOfFrame = videoIn_fork_io_outputs_0_payload_frame_endOfFrame;
  assign in2fifoAdded_payload_endOfPack = videoIn_fork_io_outputs_0_payload_endOfPack;
  always @(*) begin
    fifo2outThrown_valid = fifo_pop_fork_io_outputs_1_valid;
    if(fifo2outThrowCond) begin
      fifo2outThrown_valid = 1'b0;
    end
  end

  always @(*) begin
    fifo_pop_fork_io_outputs_1_ready = fifo2outThrown_ready;
    if(fifo2outThrowCond) begin
      fifo_pop_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign fifo2outThrown_payload_0_pixel_0 = fifo_pop_fork_io_outputs_1_payload_0_pixel_0;
  assign fifo2outThrown_payload_0_pixel_1 = fifo_pop_fork_io_outputs_1_payload_0_pixel_1;
  assign fifo2outThrown_payload_0_pixel_2 = fifo_pop_fork_io_outputs_1_payload_0_pixel_2;
  assign fifo2outThrown_payload_0_pixel_3 = fifo_pop_fork_io_outputs_1_payload_0_pixel_3;
  assign fifo2outThrown_payload_0_pixel_4 = fifo_pop_fork_io_outputs_1_payload_0_pixel_4;
  assign fifo2outThrown_payload_0_pixel_5 = fifo_pop_fork_io_outputs_1_payload_0_pixel_5;
  assign fifo2outThrown_payload_0_pixel_6 = fifo_pop_fork_io_outputs_1_payload_0_pixel_6;
  assign fifo2outThrown_payload_0_pixel_7 = fifo_pop_fork_io_outputs_1_payload_0_pixel_7;
  assign fifo2outThrown_payload_0_pixel_8 = fifo_pop_fork_io_outputs_1_payload_0_pixel_8;
  assign fifo2outThrown_payload_0_pixel_9 = fifo_pop_fork_io_outputs_1_payload_0_pixel_9;
  assign fifo2outThrown_payload_0_pixel_10 = fifo_pop_fork_io_outputs_1_payload_0_pixel_10;
  assign fifo2outThrown_payload_0_pixel_11 = fifo_pop_fork_io_outputs_1_payload_0_pixel_11;
  assign fifo2outThrown_payload_0_pixel_12 = fifo_pop_fork_io_outputs_1_payload_0_pixel_12;
  assign fifo2outThrown_payload_0_pixel_13 = fifo_pop_fork_io_outputs_1_payload_0_pixel_13;
  assign fifo2outThrown_payload_0_pixel_14 = fifo_pop_fork_io_outputs_1_payload_0_pixel_14;
  assign fifo2outThrown_payload_0_pixel_15 = fifo_pop_fork_io_outputs_1_payload_0_pixel_15;
  assign fifo2outThrown_payload_0_endOfLine = fifo_pop_fork_io_outputs_1_payload_0_endOfLine;
  assign fifo2outThrown_payload_1_pixel_0 = fifo_pop_fork_io_outputs_1_payload_1_pixel_0;
  assign fifo2outThrown_payload_1_pixel_1 = fifo_pop_fork_io_outputs_1_payload_1_pixel_1;
  assign fifo2outThrown_payload_1_pixel_2 = fifo_pop_fork_io_outputs_1_payload_1_pixel_2;
  assign fifo2outThrown_payload_1_pixel_3 = fifo_pop_fork_io_outputs_1_payload_1_pixel_3;
  assign fifo2outThrown_payload_1_pixel_4 = fifo_pop_fork_io_outputs_1_payload_1_pixel_4;
  assign fifo2outThrown_payload_1_pixel_5 = fifo_pop_fork_io_outputs_1_payload_1_pixel_5;
  assign fifo2outThrown_payload_1_pixel_6 = fifo_pop_fork_io_outputs_1_payload_1_pixel_6;
  assign fifo2outThrown_payload_1_pixel_7 = fifo_pop_fork_io_outputs_1_payload_1_pixel_7;
  assign fifo2outThrown_payload_1_pixel_8 = fifo_pop_fork_io_outputs_1_payload_1_pixel_8;
  assign fifo2outThrown_payload_1_pixel_9 = fifo_pop_fork_io_outputs_1_payload_1_pixel_9;
  assign fifo2outThrown_payload_1_pixel_10 = fifo_pop_fork_io_outputs_1_payload_1_pixel_10;
  assign fifo2outThrown_payload_1_pixel_11 = fifo_pop_fork_io_outputs_1_payload_1_pixel_11;
  assign fifo2outThrown_payload_1_pixel_12 = fifo_pop_fork_io_outputs_1_payload_1_pixel_12;
  assign fifo2outThrown_payload_1_pixel_13 = fifo_pop_fork_io_outputs_1_payload_1_pixel_13;
  assign fifo2outThrown_payload_1_pixel_14 = fifo_pop_fork_io_outputs_1_payload_1_pixel_14;
  assign fifo2outThrown_payload_1_pixel_15 = fifo_pop_fork_io_outputs_1_payload_1_pixel_15;
  assign fifo2outThrown_payload_1_endOfLine = fifo_pop_fork_io_outputs_1_payload_1_endOfLine;
  always @(*) begin
    tmp_feedbackThrownAdded_valid = fifo_pop_fork_io_outputs_0_valid;
    if(feedbackThrowCond) begin
      tmp_feedbackThrownAdded_valid = 1'b0;
    end
  end

  always @(*) begin
    fifo_pop_fork_io_outputs_0_ready = tmp_io_outputs_0_ready;
    if(feedbackThrowCond) begin
      fifo_pop_fork_io_outputs_0_ready = 1'b1;
    end
  end

  always @(*) begin
    feedbackThrownAdded_valid = tmp_feedbackThrownAdded_valid;
    if(feedbackAddCond) begin
      feedbackThrownAdded_valid = 1'b1;
    end
  end

  always @(*) begin
    tmp_io_outputs_0_ready = feedbackThrownAdded_ready;
    if(feedbackAddCond) begin
      tmp_io_outputs_0_ready = 1'b0;
    end
  end

  assign feedbackThrownAdded_payload_0_pixel_0 = fifo_pop_fork_io_outputs_0_payload_0_pixel_0;
  assign feedbackThrownAdded_payload_0_pixel_1 = fifo_pop_fork_io_outputs_0_payload_0_pixel_1;
  assign feedbackThrownAdded_payload_0_pixel_2 = fifo_pop_fork_io_outputs_0_payload_0_pixel_2;
  assign feedbackThrownAdded_payload_0_pixel_3 = fifo_pop_fork_io_outputs_0_payload_0_pixel_3;
  assign feedbackThrownAdded_payload_0_pixel_4 = fifo_pop_fork_io_outputs_0_payload_0_pixel_4;
  assign feedbackThrownAdded_payload_0_pixel_5 = fifo_pop_fork_io_outputs_0_payload_0_pixel_5;
  assign feedbackThrownAdded_payload_0_pixel_6 = fifo_pop_fork_io_outputs_0_payload_0_pixel_6;
  assign feedbackThrownAdded_payload_0_pixel_7 = fifo_pop_fork_io_outputs_0_payload_0_pixel_7;
  assign feedbackThrownAdded_payload_0_pixel_8 = fifo_pop_fork_io_outputs_0_payload_0_pixel_8;
  assign feedbackThrownAdded_payload_0_pixel_9 = fifo_pop_fork_io_outputs_0_payload_0_pixel_9;
  assign feedbackThrownAdded_payload_0_pixel_10 = fifo_pop_fork_io_outputs_0_payload_0_pixel_10;
  assign feedbackThrownAdded_payload_0_pixel_11 = fifo_pop_fork_io_outputs_0_payload_0_pixel_11;
  assign feedbackThrownAdded_payload_0_pixel_12 = fifo_pop_fork_io_outputs_0_payload_0_pixel_12;
  assign feedbackThrownAdded_payload_0_pixel_13 = fifo_pop_fork_io_outputs_0_payload_0_pixel_13;
  assign feedbackThrownAdded_payload_0_pixel_14 = fifo_pop_fork_io_outputs_0_payload_0_pixel_14;
  assign feedbackThrownAdded_payload_0_pixel_15 = fifo_pop_fork_io_outputs_0_payload_0_pixel_15;
  assign feedbackThrownAdded_payload_0_endOfLine = fifo_pop_fork_io_outputs_0_payload_0_endOfLine;
  assign feedbackThrownAdded_payload_1_pixel_0 = fifo_pop_fork_io_outputs_0_payload_1_pixel_0;
  assign feedbackThrownAdded_payload_1_pixel_1 = fifo_pop_fork_io_outputs_0_payload_1_pixel_1;
  assign feedbackThrownAdded_payload_1_pixel_2 = fifo_pop_fork_io_outputs_0_payload_1_pixel_2;
  assign feedbackThrownAdded_payload_1_pixel_3 = fifo_pop_fork_io_outputs_0_payload_1_pixel_3;
  assign feedbackThrownAdded_payload_1_pixel_4 = fifo_pop_fork_io_outputs_0_payload_1_pixel_4;
  assign feedbackThrownAdded_payload_1_pixel_5 = fifo_pop_fork_io_outputs_0_payload_1_pixel_5;
  assign feedbackThrownAdded_payload_1_pixel_6 = fifo_pop_fork_io_outputs_0_payload_1_pixel_6;
  assign feedbackThrownAdded_payload_1_pixel_7 = fifo_pop_fork_io_outputs_0_payload_1_pixel_7;
  assign feedbackThrownAdded_payload_1_pixel_8 = fifo_pop_fork_io_outputs_0_payload_1_pixel_8;
  assign feedbackThrownAdded_payload_1_pixel_9 = fifo_pop_fork_io_outputs_0_payload_1_pixel_9;
  assign feedbackThrownAdded_payload_1_pixel_10 = fifo_pop_fork_io_outputs_0_payload_1_pixel_10;
  assign feedbackThrownAdded_payload_1_pixel_11 = fifo_pop_fork_io_outputs_0_payload_1_pixel_11;
  assign feedbackThrownAdded_payload_1_pixel_12 = fifo_pop_fork_io_outputs_0_payload_1_pixel_12;
  assign feedbackThrownAdded_payload_1_pixel_13 = fifo_pop_fork_io_outputs_0_payload_1_pixel_13;
  assign feedbackThrownAdded_payload_1_pixel_14 = fifo_pop_fork_io_outputs_0_payload_1_pixel_14;
  assign feedbackThrownAdded_payload_1_pixel_15 = fifo_pop_fork_io_outputs_0_payload_1_pixel_15;
  assign feedbackThrownAdded_payload_1_endOfLine = fifo_pop_fork_io_outputs_0_payload_1_endOfLine;
  assign in2fifoJoinFeedback_valid = (in2fifoAdded_valid && feedbackThrownAdded_valid);
  assign in2fifoJoinFeedback_fire = (in2fifoJoinFeedback_valid && in2fifoJoinFeedback_ready);
  assign in2fifoAdded_ready = in2fifoJoinFeedback_fire;
  assign in2fifoJoinFeedback_fire_1 = (in2fifoJoinFeedback_valid && in2fifoJoinFeedback_ready);
  assign feedbackThrownAdded_ready = in2fifoJoinFeedback_fire_1;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_0 = in2fifoAdded_payload_frame_line_pixel_0;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_1 = in2fifoAdded_payload_frame_line_pixel_1;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_2 = in2fifoAdded_payload_frame_line_pixel_2;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_3 = in2fifoAdded_payload_frame_line_pixel_3;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_4 = in2fifoAdded_payload_frame_line_pixel_4;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_5 = in2fifoAdded_payload_frame_line_pixel_5;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_6 = in2fifoAdded_payload_frame_line_pixel_6;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_7 = in2fifoAdded_payload_frame_line_pixel_7;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_8 = in2fifoAdded_payload_frame_line_pixel_8;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_9 = in2fifoAdded_payload_frame_line_pixel_9;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_10 = in2fifoAdded_payload_frame_line_pixel_10;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_11 = in2fifoAdded_payload_frame_line_pixel_11;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_12 = in2fifoAdded_payload_frame_line_pixel_12;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_13 = in2fifoAdded_payload_frame_line_pixel_13;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_14 = in2fifoAdded_payload_frame_line_pixel_14;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_15 = in2fifoAdded_payload_frame_line_pixel_15;
  assign in2fifoJoinFeedback_payload__1_frame_line_endOfLine = in2fifoAdded_payload_frame_line_endOfLine;
  assign in2fifoJoinFeedback_payload__1_frame_endOfFrame = in2fifoAdded_payload_frame_endOfFrame;
  assign in2fifoJoinFeedback_payload__1_endOfPack = in2fifoAdded_payload_endOfPack;
  assign in2fifoJoinFeedback_payload__2_0_pixel_0 = feedbackThrownAdded_payload_0_pixel_0;
  assign in2fifoJoinFeedback_payload__2_0_pixel_1 = feedbackThrownAdded_payload_0_pixel_1;
  assign in2fifoJoinFeedback_payload__2_0_pixel_2 = feedbackThrownAdded_payload_0_pixel_2;
  assign in2fifoJoinFeedback_payload__2_0_pixel_3 = feedbackThrownAdded_payload_0_pixel_3;
  assign in2fifoJoinFeedback_payload__2_0_pixel_4 = feedbackThrownAdded_payload_0_pixel_4;
  assign in2fifoJoinFeedback_payload__2_0_pixel_5 = feedbackThrownAdded_payload_0_pixel_5;
  assign in2fifoJoinFeedback_payload__2_0_pixel_6 = feedbackThrownAdded_payload_0_pixel_6;
  assign in2fifoJoinFeedback_payload__2_0_pixel_7 = feedbackThrownAdded_payload_0_pixel_7;
  assign in2fifoJoinFeedback_payload__2_0_pixel_8 = feedbackThrownAdded_payload_0_pixel_8;
  assign in2fifoJoinFeedback_payload__2_0_pixel_9 = feedbackThrownAdded_payload_0_pixel_9;
  assign in2fifoJoinFeedback_payload__2_0_pixel_10 = feedbackThrownAdded_payload_0_pixel_10;
  assign in2fifoJoinFeedback_payload__2_0_pixel_11 = feedbackThrownAdded_payload_0_pixel_11;
  assign in2fifoJoinFeedback_payload__2_0_pixel_12 = feedbackThrownAdded_payload_0_pixel_12;
  assign in2fifoJoinFeedback_payload__2_0_pixel_13 = feedbackThrownAdded_payload_0_pixel_13;
  assign in2fifoJoinFeedback_payload__2_0_pixel_14 = feedbackThrownAdded_payload_0_pixel_14;
  assign in2fifoJoinFeedback_payload__2_0_pixel_15 = feedbackThrownAdded_payload_0_pixel_15;
  assign in2fifoJoinFeedback_payload__2_0_endOfLine = feedbackThrownAdded_payload_0_endOfLine;
  assign in2fifoJoinFeedback_payload__2_1_pixel_0 = feedbackThrownAdded_payload_1_pixel_0;
  assign in2fifoJoinFeedback_payload__2_1_pixel_1 = feedbackThrownAdded_payload_1_pixel_1;
  assign in2fifoJoinFeedback_payload__2_1_pixel_2 = feedbackThrownAdded_payload_1_pixel_2;
  assign in2fifoJoinFeedback_payload__2_1_pixel_3 = feedbackThrownAdded_payload_1_pixel_3;
  assign in2fifoJoinFeedback_payload__2_1_pixel_4 = feedbackThrownAdded_payload_1_pixel_4;
  assign in2fifoJoinFeedback_payload__2_1_pixel_5 = feedbackThrownAdded_payload_1_pixel_5;
  assign in2fifoJoinFeedback_payload__2_1_pixel_6 = feedbackThrownAdded_payload_1_pixel_6;
  assign in2fifoJoinFeedback_payload__2_1_pixel_7 = feedbackThrownAdded_payload_1_pixel_7;
  assign in2fifoJoinFeedback_payload__2_1_pixel_8 = feedbackThrownAdded_payload_1_pixel_8;
  assign in2fifoJoinFeedback_payload__2_1_pixel_9 = feedbackThrownAdded_payload_1_pixel_9;
  assign in2fifoJoinFeedback_payload__2_1_pixel_10 = feedbackThrownAdded_payload_1_pixel_10;
  assign in2fifoJoinFeedback_payload__2_1_pixel_11 = feedbackThrownAdded_payload_1_pixel_11;
  assign in2fifoJoinFeedback_payload__2_1_pixel_12 = feedbackThrownAdded_payload_1_pixel_12;
  assign in2fifoJoinFeedback_payload__2_1_pixel_13 = feedbackThrownAdded_payload_1_pixel_13;
  assign in2fifoJoinFeedback_payload__2_1_pixel_14 = feedbackThrownAdded_payload_1_pixel_14;
  assign in2fifoJoinFeedback_payload__2_1_pixel_15 = feedbackThrownAdded_payload_1_pixel_15;
  assign in2fifoJoinFeedback_payload__2_1_endOfLine = feedbackThrownAdded_payload_1_endOfLine;
  assign in2outJoinFifo2out_valid = (in2outThrownAdded_valid && fifo2outThrown_valid);
  assign in2outJoinFifo2out_fire = (in2outJoinFifo2out_valid && in2outJoinFifo2out_ready);
  assign in2outThrownAdded_ready = in2outJoinFifo2out_fire;
  assign in2outJoinFifo2out_fire_1 = (in2outJoinFifo2out_valid && in2outJoinFifo2out_ready);
  assign fifo2outThrown_ready = in2outJoinFifo2out_fire_1;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_0 = in2outThrownAdded_payload_frame_line_pixel_0;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_1 = in2outThrownAdded_payload_frame_line_pixel_1;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_2 = in2outThrownAdded_payload_frame_line_pixel_2;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_3 = in2outThrownAdded_payload_frame_line_pixel_3;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_4 = in2outThrownAdded_payload_frame_line_pixel_4;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_5 = in2outThrownAdded_payload_frame_line_pixel_5;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_6 = in2outThrownAdded_payload_frame_line_pixel_6;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_7 = in2outThrownAdded_payload_frame_line_pixel_7;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_8 = in2outThrownAdded_payload_frame_line_pixel_8;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_9 = in2outThrownAdded_payload_frame_line_pixel_9;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_10 = in2outThrownAdded_payload_frame_line_pixel_10;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_11 = in2outThrownAdded_payload_frame_line_pixel_11;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_12 = in2outThrownAdded_payload_frame_line_pixel_12;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_13 = in2outThrownAdded_payload_frame_line_pixel_13;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_14 = in2outThrownAdded_payload_frame_line_pixel_14;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_15 = in2outThrownAdded_payload_frame_line_pixel_15;
  assign in2outJoinFifo2out_payload__1_frame_line_endOfLine = in2outThrownAdded_payload_frame_line_endOfLine;
  assign in2outJoinFifo2out_payload__1_frame_endOfFrame = in2outThrownAdded_payload_frame_endOfFrame;
  assign in2outJoinFifo2out_payload__1_endOfPack = in2outThrownAdded_payload_endOfPack;
  assign in2outJoinFifo2out_payload__2_0_pixel_0 = fifo2outThrown_payload_0_pixel_0;
  assign in2outJoinFifo2out_payload__2_0_pixel_1 = fifo2outThrown_payload_0_pixel_1;
  assign in2outJoinFifo2out_payload__2_0_pixel_2 = fifo2outThrown_payload_0_pixel_2;
  assign in2outJoinFifo2out_payload__2_0_pixel_3 = fifo2outThrown_payload_0_pixel_3;
  assign in2outJoinFifo2out_payload__2_0_pixel_4 = fifo2outThrown_payload_0_pixel_4;
  assign in2outJoinFifo2out_payload__2_0_pixel_5 = fifo2outThrown_payload_0_pixel_5;
  assign in2outJoinFifo2out_payload__2_0_pixel_6 = fifo2outThrown_payload_0_pixel_6;
  assign in2outJoinFifo2out_payload__2_0_pixel_7 = fifo2outThrown_payload_0_pixel_7;
  assign in2outJoinFifo2out_payload__2_0_pixel_8 = fifo2outThrown_payload_0_pixel_8;
  assign in2outJoinFifo2out_payload__2_0_pixel_9 = fifo2outThrown_payload_0_pixel_9;
  assign in2outJoinFifo2out_payload__2_0_pixel_10 = fifo2outThrown_payload_0_pixel_10;
  assign in2outJoinFifo2out_payload__2_0_pixel_11 = fifo2outThrown_payload_0_pixel_11;
  assign in2outJoinFifo2out_payload__2_0_pixel_12 = fifo2outThrown_payload_0_pixel_12;
  assign in2outJoinFifo2out_payload__2_0_pixel_13 = fifo2outThrown_payload_0_pixel_13;
  assign in2outJoinFifo2out_payload__2_0_pixel_14 = fifo2outThrown_payload_0_pixel_14;
  assign in2outJoinFifo2out_payload__2_0_pixel_15 = fifo2outThrown_payload_0_pixel_15;
  assign in2outJoinFifo2out_payload__2_0_endOfLine = fifo2outThrown_payload_0_endOfLine;
  assign in2outJoinFifo2out_payload__2_1_pixel_0 = fifo2outThrown_payload_1_pixel_0;
  assign in2outJoinFifo2out_payload__2_1_pixel_1 = fifo2outThrown_payload_1_pixel_1;
  assign in2outJoinFifo2out_payload__2_1_pixel_2 = fifo2outThrown_payload_1_pixel_2;
  assign in2outJoinFifo2out_payload__2_1_pixel_3 = fifo2outThrown_payload_1_pixel_3;
  assign in2outJoinFifo2out_payload__2_1_pixel_4 = fifo2outThrown_payload_1_pixel_4;
  assign in2outJoinFifo2out_payload__2_1_pixel_5 = fifo2outThrown_payload_1_pixel_5;
  assign in2outJoinFifo2out_payload__2_1_pixel_6 = fifo2outThrown_payload_1_pixel_6;
  assign in2outJoinFifo2out_payload__2_1_pixel_7 = fifo2outThrown_payload_1_pixel_7;
  assign in2outJoinFifo2out_payload__2_1_pixel_8 = fifo2outThrown_payload_1_pixel_8;
  assign in2outJoinFifo2out_payload__2_1_pixel_9 = fifo2outThrown_payload_1_pixel_9;
  assign in2outJoinFifo2out_payload__2_1_pixel_10 = fifo2outThrown_payload_1_pixel_10;
  assign in2outJoinFifo2out_payload__2_1_pixel_11 = fifo2outThrown_payload_1_pixel_11;
  assign in2outJoinFifo2out_payload__2_1_pixel_12 = fifo2outThrown_payload_1_pixel_12;
  assign in2outJoinFifo2out_payload__2_1_pixel_13 = fifo2outThrown_payload_1_pixel_13;
  assign in2outJoinFifo2out_payload__2_1_pixel_14 = fifo2outThrown_payload_1_pixel_14;
  assign in2outJoinFifo2out_payload__2_1_pixel_15 = fifo2outThrown_payload_1_pixel_15;
  assign in2outJoinFifo2out_payload__2_1_endOfLine = fifo2outThrown_payload_1_endOfLine;
  always @(*) begin
    firstFewLines_willIncrement = 1'b0;
    if(when_LineBufferSame_l72) begin
      firstFewLines_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    firstFewLines_willClear = 1'b0;
    if(when_LineBufferSame_l71) begin
      firstFewLines_willClear = 1'b1;
    end
  end

  assign firstFewLines_willOverflowIfInc = (firstFewLines_value == 1'b1);
  assign firstFewLines_willOverflow = (firstFewLines_willOverflowIfInc && firstFewLines_willIncrement);
  always @(*) begin
    firstFewLines_valueNext = (firstFewLines_value + firstFewLines_willIncrement);
    if(firstFewLines_willClear) begin
      firstFewLines_valueNext = 1'b0;
    end
  end

  assign ioVideoInFire = (videoIn_valid && videoIn_ready);
  assign firstLine = (firstFewLines_value == 1'b0);
  assign firstFewLinesWontOverflowIfInc = (! firstFewLines_willOverflowIfInc);
  assign when_LineBufferSame_l71 = (ioVideoInFire && videoIn_payload_endOfPack);
  assign when_LineBufferSame_l72 = ((ioVideoInFire && videoIn_payload_frame_line_endOfLine) && firstFewLinesWontOverflowIfInc);
  always @(*) begin
    lastFewLines_willIncrement = 1'b0;
    if(when_LineBufferSame_l78) begin
      lastFewLines_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    lastFewLines_willClear = 1'b0;
    if(when_LineBufferSame_l77) begin
      lastFewLines_willClear = 1'b1;
    end
  end

  assign lastFewLines_willOverflowIfInc = 1'b1;
  assign lastFewLines_willOverflow = (lastFewLines_willOverflowIfInc && lastFewLines_willIncrement);
  assign ioVideoOutFire = (videoOut_valid && videoOut_ready);
  assign lastFewLinesWontOverflowIfInc = (! lastFewLines_willOverflowIfInc);
  assign when_LineBufferSame_l77 = (ioVideoOutFire && in2outJoinFifo2out_payload__1_frame_endOfFrame);
  assign when_LineBufferSame_l78 = (ioVideoOutFire && in2outJoinFifo2out_payload__2_1_endOfLine);
  assign when_LineBufferSame_l81 = (ioVideoInFire && videoIn_payload_frame_endOfFrame);
  assign when_LineBufferSame_l81_1 = (ioVideoOutFire && videoOut_payload_frame_endOfFrame);
  assign when_LineBufferSame_l83 = (ioVideoInFire && videoIn_payload_endOfPack);
  assign when_LineBufferSame_l83_1 = (ioVideoOutFire && videoOut_payload_endOfPack);
  assign endOfPackGapInv = (! endOfPackGap);
  assign in2outThrowCond = (endOfPackGapInv && firstFewLinesWontOverflowIfInc);
  assign feedbackAddCond = (endOfPackGapInv && firstLine);
  assign fifo2outThrowCond = ((endOfPackGapInv && (! firstLine)) && firstFewLinesWontOverflowIfInc);
  assign in2outAddCond = endOfPackGap;
  assign feedbackThrowCond = (endOfPackGap && lastFewLines_willOverflowIfInc);
  assign in2fifoAddCond = (endOfPackGap && lastFewLinesWontOverflowIfInc);
  assign in2fifoJoinFeedback_ready = fifo_push_ready;
  assign cntPrevStable = (cntPrev == 2'b01);
  assign cntPostStable = (cntPost == 2'b01);
  assign cntPrevEqualVec_0 = ((2'b00 <= cntPrev) && (cntPrev < 2'b01));
  assign cntPostEqualVec_0 = (cntPost <= 2'b00);
  assign when_LineBufferSame_l103 = (ioVideoInFire && videoIn_payload_frame_endOfFrame);
  assign when_LineBufferSame_l104 = (ioVideoOutFire && videoOut_payload_frame_endOfFrame);
  assign when_LineBufferSame_l105 = ((ioVideoOutFire && videoOut_payload_frame_line_endOfLine) && (! cntPrevStable));
  assign when_LineBufferSame_l106 = ((ioVideoOutFire && videoOut_payload_frame_line_endOfLine) && (! cntPostStable));
  assign up_0_0 = (cntPostEqualVec_0 ? zero_0 : in2outJoinFifo2out_payload__2_0_pixel_0);
  assign up_0_1 = (cntPostEqualVec_0 ? zero_1 : in2outJoinFifo2out_payload__2_0_pixel_1);
  assign up_0_2 = (cntPostEqualVec_0 ? zero_2 : in2outJoinFifo2out_payload__2_0_pixel_2);
  assign up_0_3 = (cntPostEqualVec_0 ? zero_3 : in2outJoinFifo2out_payload__2_0_pixel_3);
  assign up_0_4 = (cntPostEqualVec_0 ? zero_4 : in2outJoinFifo2out_payload__2_0_pixel_4);
  assign up_0_5 = (cntPostEqualVec_0 ? zero_5 : in2outJoinFifo2out_payload__2_0_pixel_5);
  assign up_0_6 = (cntPostEqualVec_0 ? zero_6 : in2outJoinFifo2out_payload__2_0_pixel_6);
  assign up_0_7 = (cntPostEqualVec_0 ? zero_7 : in2outJoinFifo2out_payload__2_0_pixel_7);
  assign up_0_8 = (cntPostEqualVec_0 ? zero_8 : in2outJoinFifo2out_payload__2_0_pixel_8);
  assign up_0_9 = (cntPostEqualVec_0 ? zero_9 : in2outJoinFifo2out_payload__2_0_pixel_9);
  assign up_0_10 = (cntPostEqualVec_0 ? zero_10 : in2outJoinFifo2out_payload__2_0_pixel_10);
  assign up_0_11 = (cntPostEqualVec_0 ? zero_11 : in2outJoinFifo2out_payload__2_0_pixel_11);
  assign up_0_12 = (cntPostEqualVec_0 ? zero_12 : in2outJoinFifo2out_payload__2_0_pixel_12);
  assign up_0_13 = (cntPostEqualVec_0 ? zero_13 : in2outJoinFifo2out_payload__2_0_pixel_13);
  assign up_0_14 = (cntPostEqualVec_0 ? zero_14 : in2outJoinFifo2out_payload__2_0_pixel_14);
  assign up_0_15 = (cntPostEqualVec_0 ? zero_15 : in2outJoinFifo2out_payload__2_0_pixel_15);
  assign down_0_0 = (cntPrevEqualVec_0 ? zero_0 : in2outJoinFifo2out_payload__1_frame_line_pixel_0);
  assign down_0_1 = (cntPrevEqualVec_0 ? zero_1 : in2outJoinFifo2out_payload__1_frame_line_pixel_1);
  assign down_0_2 = (cntPrevEqualVec_0 ? zero_2 : in2outJoinFifo2out_payload__1_frame_line_pixel_2);
  assign down_0_3 = (cntPrevEqualVec_0 ? zero_3 : in2outJoinFifo2out_payload__1_frame_line_pixel_3);
  assign down_0_4 = (cntPrevEqualVec_0 ? zero_4 : in2outJoinFifo2out_payload__1_frame_line_pixel_4);
  assign down_0_5 = (cntPrevEqualVec_0 ? zero_5 : in2outJoinFifo2out_payload__1_frame_line_pixel_5);
  assign down_0_6 = (cntPrevEqualVec_0 ? zero_6 : in2outJoinFifo2out_payload__1_frame_line_pixel_6);
  assign down_0_7 = (cntPrevEqualVec_0 ? zero_7 : in2outJoinFifo2out_payload__1_frame_line_pixel_7);
  assign down_0_8 = (cntPrevEqualVec_0 ? zero_8 : in2outJoinFifo2out_payload__1_frame_line_pixel_8);
  assign down_0_9 = (cntPrevEqualVec_0 ? zero_9 : in2outJoinFifo2out_payload__1_frame_line_pixel_9);
  assign down_0_10 = (cntPrevEqualVec_0 ? zero_10 : in2outJoinFifo2out_payload__1_frame_line_pixel_10);
  assign down_0_11 = (cntPrevEqualVec_0 ? zero_11 : in2outJoinFifo2out_payload__1_frame_line_pixel_11);
  assign down_0_12 = (cntPrevEqualVec_0 ? zero_12 : in2outJoinFifo2out_payload__1_frame_line_pixel_12);
  assign down_0_13 = (cntPrevEqualVec_0 ? zero_13 : in2outJoinFifo2out_payload__1_frame_line_pixel_13);
  assign down_0_14 = (cntPrevEqualVec_0 ? zero_14 : in2outJoinFifo2out_payload__1_frame_line_pixel_14);
  assign down_0_15 = (cntPrevEqualVec_0 ? zero_15 : in2outJoinFifo2out_payload__1_frame_line_pixel_15);
  assign videoOut_valid = in2outJoinFifo2out_valid;
  assign in2outJoinFifo2out_ready = videoOut_ready;
  assign videoOut_payload_endOfPack = ((endOfPackGap && videoOut_payload_frame_line_endOfLine) && lastFewLines_willOverflowIfInc);
  assign videoOut_payload_frame_endOfFrame = ((endOfFrameGap && videoOut_payload_frame_line_endOfLine) && lastFewLines_willOverflowIfInc);
  assign videoOut_payload_frame_line_pixel_0_0 = up_0_0;
  assign videoOut_payload_frame_line_pixel_0_1 = up_0_1;
  assign videoOut_payload_frame_line_pixel_0_2 = up_0_2;
  assign videoOut_payload_frame_line_pixel_0_3 = up_0_3;
  assign videoOut_payload_frame_line_pixel_0_4 = up_0_4;
  assign videoOut_payload_frame_line_pixel_0_5 = up_0_5;
  assign videoOut_payload_frame_line_pixel_0_6 = up_0_6;
  assign videoOut_payload_frame_line_pixel_0_7 = up_0_7;
  assign videoOut_payload_frame_line_pixel_0_8 = up_0_8;
  assign videoOut_payload_frame_line_pixel_0_9 = up_0_9;
  assign videoOut_payload_frame_line_pixel_0_10 = up_0_10;
  assign videoOut_payload_frame_line_pixel_0_11 = up_0_11;
  assign videoOut_payload_frame_line_pixel_0_12 = up_0_12;
  assign videoOut_payload_frame_line_pixel_0_13 = up_0_13;
  assign videoOut_payload_frame_line_pixel_0_14 = up_0_14;
  assign videoOut_payload_frame_line_pixel_0_15 = up_0_15;
  assign videoOut_payload_frame_line_pixel_1_0 = in2outJoinFifo2out_payload__2_1_pixel_0;
  assign videoOut_payload_frame_line_pixel_1_1 = in2outJoinFifo2out_payload__2_1_pixel_1;
  assign videoOut_payload_frame_line_pixel_1_2 = in2outJoinFifo2out_payload__2_1_pixel_2;
  assign videoOut_payload_frame_line_pixel_1_3 = in2outJoinFifo2out_payload__2_1_pixel_3;
  assign videoOut_payload_frame_line_pixel_1_4 = in2outJoinFifo2out_payload__2_1_pixel_4;
  assign videoOut_payload_frame_line_pixel_1_5 = in2outJoinFifo2out_payload__2_1_pixel_5;
  assign videoOut_payload_frame_line_pixel_1_6 = in2outJoinFifo2out_payload__2_1_pixel_6;
  assign videoOut_payload_frame_line_pixel_1_7 = in2outJoinFifo2out_payload__2_1_pixel_7;
  assign videoOut_payload_frame_line_pixel_1_8 = in2outJoinFifo2out_payload__2_1_pixel_8;
  assign videoOut_payload_frame_line_pixel_1_9 = in2outJoinFifo2out_payload__2_1_pixel_9;
  assign videoOut_payload_frame_line_pixel_1_10 = in2outJoinFifo2out_payload__2_1_pixel_10;
  assign videoOut_payload_frame_line_pixel_1_11 = in2outJoinFifo2out_payload__2_1_pixel_11;
  assign videoOut_payload_frame_line_pixel_1_12 = in2outJoinFifo2out_payload__2_1_pixel_12;
  assign videoOut_payload_frame_line_pixel_1_13 = in2outJoinFifo2out_payload__2_1_pixel_13;
  assign videoOut_payload_frame_line_pixel_1_14 = in2outJoinFifo2out_payload__2_1_pixel_14;
  assign videoOut_payload_frame_line_pixel_1_15 = in2outJoinFifo2out_payload__2_1_pixel_15;
  assign videoOut_payload_frame_line_pixel_2_0 = down_0_0;
  assign videoOut_payload_frame_line_pixel_2_1 = down_0_1;
  assign videoOut_payload_frame_line_pixel_2_2 = down_0_2;
  assign videoOut_payload_frame_line_pixel_2_3 = down_0_3;
  assign videoOut_payload_frame_line_pixel_2_4 = down_0_4;
  assign videoOut_payload_frame_line_pixel_2_5 = down_0_5;
  assign videoOut_payload_frame_line_pixel_2_6 = down_0_6;
  assign videoOut_payload_frame_line_pixel_2_7 = down_0_7;
  assign videoOut_payload_frame_line_pixel_2_8 = down_0_8;
  assign videoOut_payload_frame_line_pixel_2_9 = down_0_9;
  assign videoOut_payload_frame_line_pixel_2_10 = down_0_10;
  assign videoOut_payload_frame_line_pixel_2_11 = down_0_11;
  assign videoOut_payload_frame_line_pixel_2_12 = down_0_12;
  assign videoOut_payload_frame_line_pixel_2_13 = down_0_13;
  assign videoOut_payload_frame_line_pixel_2_14 = down_0_14;
  assign videoOut_payload_frame_line_pixel_2_15 = down_0_15;
  assign videoOut_payload_frame_line_endOfLine = in2outJoinFifo2out_payload__2_1_endOfLine;
  always @(posedge clk) begin
    if(reset) begin
      firstFewLines_value <= 1'b0;
      endOfFrameGap <= 1'b0;
      endOfPackGap <= 1'b0;
      cntPrev <= 2'b01;
      cntPost <= 2'b00;
    end else begin
      firstFewLines_value <= firstFewLines_valueNext;
      if(when_LineBufferSame_l81) begin
        endOfFrameGap <= 1'b1;
      end
      if(when_LineBufferSame_l81_1) begin
        endOfFrameGap <= 1'b0;
      end
      if(when_LineBufferSame_l83) begin
        endOfPackGap <= 1'b1;
      end
      if(when_LineBufferSame_l83_1) begin
        endOfPackGap <= 1'b0;
      end
      if(when_LineBufferSame_l103) begin
        cntPrev <= 2'b00;
      end
      if(when_LineBufferSame_l104) begin
        cntPost <= 2'b00;
      end
      if(when_LineBufferSame_l105) begin
        cntPrev <= (cntPrev + 2'b01);
      end
      if(when_LineBufferSame_l106) begin
        cntPost <= (cntPost + 2'b01);
      end
    end
  end


endmodule

module PixelBufferValid (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_0_15,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_1_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  wire       [7:0]    tmp_pixelBuffer;
  wire       [63:0]   tmp_pixelBuffer_1;
  wire       [7:0]    tmp_pixelBuffer_2;
  wire       [63:0]   tmp_pixelBuffer_3;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0;
  wire       [71:0]   tmp_tmp_pixelVec_0_0_0_1;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_2;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_3;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_4;
  wire       [71:0]   tmp_tmp_pixelVec_0_0_0_5;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_6;
  wire       [7:0]    tmp_tmp_pixelVec_0_0_0_7;
  wire                videoInFire;
  wire                videoOutFire;
  reg        [255:0]  pixelBuffer;
  wire                bridge_valid;
  reg                 bridge_ready;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    bridge_payload_frame_line_pixel_1_1_15;
  wire                bridge_payload_frame_line_endOfLine;
  wire                bridge_payload_frame_endOfFrame;
  wire                bridge_payload_endOfPack;
  wire                bridgeFire;
  reg                 pixelCnt_willIncrement;
  reg                 pixelCnt_willClear;
  reg        [0:0]    pixelCnt_valueNext;
  reg        [0:0]    pixelCnt_value;
  wire                pixelCnt_willOverflowIfInc;
  wire                pixelCnt_willOverflow;
  wire                pixelCntWontOverflowIfInc;
  wire                when_PixelBufferValid_l32;
  wire                when_PixelBufferValid_l33;
  wire       [7:0]    pixelVec_0_0_0;
  wire       [7:0]    pixelVec_0_0_1;
  wire       [7:0]    pixelVec_0_0_2;
  wire       [7:0]    pixelVec_0_0_3;
  wire       [7:0]    pixelVec_0_0_4;
  wire       [7:0]    pixelVec_0_0_5;
  wire       [7:0]    pixelVec_0_0_6;
  wire       [7:0]    pixelVec_0_0_7;
  wire       [7:0]    pixelVec_0_0_8;
  wire       [7:0]    pixelVec_0_0_9;
  wire       [7:0]    pixelVec_0_0_10;
  wire       [7:0]    pixelVec_0_0_11;
  wire       [7:0]    pixelVec_0_0_12;
  wire       [7:0]    pixelVec_0_0_13;
  wire       [7:0]    pixelVec_0_0_14;
  wire       [7:0]    pixelVec_0_0_15;
  wire       [7:0]    pixelVec_0_1_0;
  wire       [7:0]    pixelVec_0_1_1;
  wire       [7:0]    pixelVec_0_1_2;
  wire       [7:0]    pixelVec_0_1_3;
  wire       [7:0]    pixelVec_0_1_4;
  wire       [7:0]    pixelVec_0_1_5;
  wire       [7:0]    pixelVec_0_1_6;
  wire       [7:0]    pixelVec_0_1_7;
  wire       [7:0]    pixelVec_0_1_8;
  wire       [7:0]    pixelVec_0_1_9;
  wire       [7:0]    pixelVec_0_1_10;
  wire       [7:0]    pixelVec_0_1_11;
  wire       [7:0]    pixelVec_0_1_12;
  wire       [7:0]    pixelVec_0_1_13;
  wire       [7:0]    pixelVec_0_1_14;
  wire       [7:0]    pixelVec_0_1_15;
  wire       [7:0]    pixelVec_1_0_0;
  wire       [7:0]    pixelVec_1_0_1;
  wire       [7:0]    pixelVec_1_0_2;
  wire       [7:0]    pixelVec_1_0_3;
  wire       [7:0]    pixelVec_1_0_4;
  wire       [7:0]    pixelVec_1_0_5;
  wire       [7:0]    pixelVec_1_0_6;
  wire       [7:0]    pixelVec_1_0_7;
  wire       [7:0]    pixelVec_1_0_8;
  wire       [7:0]    pixelVec_1_0_9;
  wire       [7:0]    pixelVec_1_0_10;
  wire       [7:0]    pixelVec_1_0_11;
  wire       [7:0]    pixelVec_1_0_12;
  wire       [7:0]    pixelVec_1_0_13;
  wire       [7:0]    pixelVec_1_0_14;
  wire       [7:0]    pixelVec_1_0_15;
  wire       [7:0]    pixelVec_1_1_0;
  wire       [7:0]    pixelVec_1_1_1;
  wire       [7:0]    pixelVec_1_1_2;
  wire       [7:0]    pixelVec_1_1_3;
  wire       [7:0]    pixelVec_1_1_4;
  wire       [7:0]    pixelVec_1_1_5;
  wire       [7:0]    pixelVec_1_1_6;
  wire       [7:0]    pixelVec_1_1_7;
  wire       [7:0]    pixelVec_1_1_8;
  wire       [7:0]    pixelVec_1_1_9;
  wire       [7:0]    pixelVec_1_1_10;
  wire       [7:0]    pixelVec_1_1_11;
  wire       [7:0]    pixelVec_1_1_12;
  wire       [7:0]    pixelVec_1_1_13;
  wire       [7:0]    pixelVec_1_1_14;
  wire       [7:0]    pixelVec_1_1_15;
  wire       [511:0]  tmp_pixelVec_0_0_0;
  wire       [255:0]  tmp_pixelVec_0_0_0_1;
  wire       [127:0]  tmp_pixelVec_0_0_0_2;
  wire       [127:0]  tmp_pixelVec_0_1_0;
  wire       [255:0]  tmp_pixelVec_1_0_0;
  wire       [127:0]  tmp_pixelVec_1_0_0_1;
  wire       [127:0]  tmp_pixelVec_1_1_0;
  reg                 bridge_thrown_valid;
  wire                bridge_thrown_ready;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_0;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_1;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_2;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_3;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_4;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_5;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_6;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_7;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_8;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_9;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_10;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_11;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_12;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_13;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_14;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_0_15;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_0;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_1;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_2;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_3;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_4;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_5;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_6;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_7;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_8;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_9;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_10;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_11;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_12;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_13;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_14;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_0_1_15;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_0;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_1;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_2;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_3;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_4;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_5;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_6;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_7;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_8;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_9;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_10;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_11;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_12;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_13;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_14;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_0_15;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_0;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_1;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_2;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_3;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_4;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_5;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_6;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_7;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_8;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_9;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_10;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_11;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_12;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_13;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_14;
  wire       [7:0]    bridge_thrown_payload_frame_line_pixel_1_1_15;
  wire                bridge_thrown_payload_frame_line_endOfLine;
  wire                bridge_thrown_payload_frame_endOfFrame;
  wire                bridge_thrown_payload_endOfPack;

  assign tmp_pixelBuffer = videoIn_payload_frame_line_pixel_1_8;
  assign tmp_pixelBuffer_1 = {videoIn_payload_frame_line_pixel_1_7,{videoIn_payload_frame_line_pixel_1_6,{videoIn_payload_frame_line_pixel_1_5,{videoIn_payload_frame_line_pixel_1_4,{videoIn_payload_frame_line_pixel_1_3,{videoIn_payload_frame_line_pixel_1_2,{videoIn_payload_frame_line_pixel_1_1,videoIn_payload_frame_line_pixel_1_0}}}}}}};
  assign tmp_pixelBuffer_2 = videoIn_payload_frame_line_pixel_0_8;
  assign tmp_pixelBuffer_3 = {videoIn_payload_frame_line_pixel_0_7,{videoIn_payload_frame_line_pixel_0_6,{videoIn_payload_frame_line_pixel_0_5,{videoIn_payload_frame_line_pixel_0_4,{videoIn_payload_frame_line_pixel_0_3,{videoIn_payload_frame_line_pixel_0_2,{videoIn_payload_frame_line_pixel_0_1,videoIn_payload_frame_line_pixel_0_0}}}}}}};
  assign tmp_tmp_pixelVec_0_0_0 = videoIn_payload_frame_line_pixel_1_9;
  assign tmp_tmp_pixelVec_0_0_0_1 = {videoIn_payload_frame_line_pixel_1_8,{videoIn_payload_frame_line_pixel_1_7,{videoIn_payload_frame_line_pixel_1_6,{videoIn_payload_frame_line_pixel_1_5,{videoIn_payload_frame_line_pixel_1_4,{videoIn_payload_frame_line_pixel_1_3,{videoIn_payload_frame_line_pixel_1_2,{tmp_tmp_pixelVec_0_0_0_2,tmp_tmp_pixelVec_0_0_0_3}}}}}}}};
  assign tmp_tmp_pixelVec_0_0_0_4 = videoIn_payload_frame_line_pixel_0_9;
  assign tmp_tmp_pixelVec_0_0_0_5 = {videoIn_payload_frame_line_pixel_0_8,{videoIn_payload_frame_line_pixel_0_7,{videoIn_payload_frame_line_pixel_0_6,{videoIn_payload_frame_line_pixel_0_5,{videoIn_payload_frame_line_pixel_0_4,{videoIn_payload_frame_line_pixel_0_3,{videoIn_payload_frame_line_pixel_0_2,{tmp_tmp_pixelVec_0_0_0_6,tmp_tmp_pixelVec_0_0_0_7}}}}}}}};
  assign tmp_tmp_pixelVec_0_0_0_2 = videoIn_payload_frame_line_pixel_1_1;
  assign tmp_tmp_pixelVec_0_0_0_3 = videoIn_payload_frame_line_pixel_1_0;
  assign tmp_tmp_pixelVec_0_0_0_6 = videoIn_payload_frame_line_pixel_0_1;
  assign tmp_tmp_pixelVec_0_0_0_7 = videoIn_payload_frame_line_pixel_0_0;
  assign videoInFire = (videoIn_valid && videoIn_ready);
  assign videoOutFire = (videoOut_valid && videoOut_ready);
  assign bridgeFire = (bridge_valid && bridge_ready);
  assign bridge_valid = videoIn_valid;
  assign videoIn_ready = bridge_ready;
  always @(*) begin
    pixelCnt_willIncrement = 1'b0;
    if(when_PixelBufferValid_l33) begin
      pixelCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pixelCnt_willClear = 1'b0;
    if(when_PixelBufferValid_l32) begin
      pixelCnt_willClear = 1'b1;
    end
  end

  assign pixelCnt_willOverflowIfInc = (pixelCnt_value == 1'b1);
  assign pixelCnt_willOverflow = (pixelCnt_willOverflowIfInc && pixelCnt_willIncrement);
  always @(*) begin
    pixelCnt_valueNext = (pixelCnt_value + pixelCnt_willIncrement);
    if(pixelCnt_willClear) begin
      pixelCnt_valueNext = 1'b0;
    end
  end

  assign pixelCntWontOverflowIfInc = (! pixelCnt_willOverflowIfInc);
  assign when_PixelBufferValid_l32 = (videoInFire && videoIn_payload_frame_line_endOfLine);
  assign when_PixelBufferValid_l33 = (videoInFire && pixelCntWontOverflowIfInc);
  assign tmp_pixelVec_0_0_0 = {{{videoIn_payload_frame_line_pixel_1_15,{videoIn_payload_frame_line_pixel_1_14,{videoIn_payload_frame_line_pixel_1_13,{videoIn_payload_frame_line_pixel_1_12,{videoIn_payload_frame_line_pixel_1_11,{videoIn_payload_frame_line_pixel_1_10,{tmp_tmp_pixelVec_0_0_0,tmp_tmp_pixelVec_0_0_0_1}}}}}}},{videoIn_payload_frame_line_pixel_0_15,{videoIn_payload_frame_line_pixel_0_14,{videoIn_payload_frame_line_pixel_0_13,{videoIn_payload_frame_line_pixel_0_12,{videoIn_payload_frame_line_pixel_0_11,{videoIn_payload_frame_line_pixel_0_10,{tmp_tmp_pixelVec_0_0_0_4,tmp_tmp_pixelVec_0_0_0_5}}}}}}}},pixelBuffer};
  assign tmp_pixelVec_0_0_0_1 = tmp_pixelVec_0_0_0[255 : 0];
  assign tmp_pixelVec_0_0_0_2 = tmp_pixelVec_0_0_0_1[127 : 0];
  assign pixelVec_0_0_0 = tmp_pixelVec_0_0_0_2[7 : 0];
  assign pixelVec_0_0_1 = tmp_pixelVec_0_0_0_2[15 : 8];
  assign pixelVec_0_0_2 = tmp_pixelVec_0_0_0_2[23 : 16];
  assign pixelVec_0_0_3 = tmp_pixelVec_0_0_0_2[31 : 24];
  assign pixelVec_0_0_4 = tmp_pixelVec_0_0_0_2[39 : 32];
  assign pixelVec_0_0_5 = tmp_pixelVec_0_0_0_2[47 : 40];
  assign pixelVec_0_0_6 = tmp_pixelVec_0_0_0_2[55 : 48];
  assign pixelVec_0_0_7 = tmp_pixelVec_0_0_0_2[63 : 56];
  assign pixelVec_0_0_8 = tmp_pixelVec_0_0_0_2[71 : 64];
  assign pixelVec_0_0_9 = tmp_pixelVec_0_0_0_2[79 : 72];
  assign pixelVec_0_0_10 = tmp_pixelVec_0_0_0_2[87 : 80];
  assign pixelVec_0_0_11 = tmp_pixelVec_0_0_0_2[95 : 88];
  assign pixelVec_0_0_12 = tmp_pixelVec_0_0_0_2[103 : 96];
  assign pixelVec_0_0_13 = tmp_pixelVec_0_0_0_2[111 : 104];
  assign pixelVec_0_0_14 = tmp_pixelVec_0_0_0_2[119 : 112];
  assign pixelVec_0_0_15 = tmp_pixelVec_0_0_0_2[127 : 120];
  assign tmp_pixelVec_0_1_0 = tmp_pixelVec_0_0_0_1[255 : 128];
  assign pixelVec_0_1_0 = tmp_pixelVec_0_1_0[7 : 0];
  assign pixelVec_0_1_1 = tmp_pixelVec_0_1_0[15 : 8];
  assign pixelVec_0_1_2 = tmp_pixelVec_0_1_0[23 : 16];
  assign pixelVec_0_1_3 = tmp_pixelVec_0_1_0[31 : 24];
  assign pixelVec_0_1_4 = tmp_pixelVec_0_1_0[39 : 32];
  assign pixelVec_0_1_5 = tmp_pixelVec_0_1_0[47 : 40];
  assign pixelVec_0_1_6 = tmp_pixelVec_0_1_0[55 : 48];
  assign pixelVec_0_1_7 = tmp_pixelVec_0_1_0[63 : 56];
  assign pixelVec_0_1_8 = tmp_pixelVec_0_1_0[71 : 64];
  assign pixelVec_0_1_9 = tmp_pixelVec_0_1_0[79 : 72];
  assign pixelVec_0_1_10 = tmp_pixelVec_0_1_0[87 : 80];
  assign pixelVec_0_1_11 = tmp_pixelVec_0_1_0[95 : 88];
  assign pixelVec_0_1_12 = tmp_pixelVec_0_1_0[103 : 96];
  assign pixelVec_0_1_13 = tmp_pixelVec_0_1_0[111 : 104];
  assign pixelVec_0_1_14 = tmp_pixelVec_0_1_0[119 : 112];
  assign pixelVec_0_1_15 = tmp_pixelVec_0_1_0[127 : 120];
  assign tmp_pixelVec_1_0_0 = tmp_pixelVec_0_0_0[511 : 256];
  assign tmp_pixelVec_1_0_0_1 = tmp_pixelVec_1_0_0[127 : 0];
  assign pixelVec_1_0_0 = tmp_pixelVec_1_0_0_1[7 : 0];
  assign pixelVec_1_0_1 = tmp_pixelVec_1_0_0_1[15 : 8];
  assign pixelVec_1_0_2 = tmp_pixelVec_1_0_0_1[23 : 16];
  assign pixelVec_1_0_3 = tmp_pixelVec_1_0_0_1[31 : 24];
  assign pixelVec_1_0_4 = tmp_pixelVec_1_0_0_1[39 : 32];
  assign pixelVec_1_0_5 = tmp_pixelVec_1_0_0_1[47 : 40];
  assign pixelVec_1_0_6 = tmp_pixelVec_1_0_0_1[55 : 48];
  assign pixelVec_1_0_7 = tmp_pixelVec_1_0_0_1[63 : 56];
  assign pixelVec_1_0_8 = tmp_pixelVec_1_0_0_1[71 : 64];
  assign pixelVec_1_0_9 = tmp_pixelVec_1_0_0_1[79 : 72];
  assign pixelVec_1_0_10 = tmp_pixelVec_1_0_0_1[87 : 80];
  assign pixelVec_1_0_11 = tmp_pixelVec_1_0_0_1[95 : 88];
  assign pixelVec_1_0_12 = tmp_pixelVec_1_0_0_1[103 : 96];
  assign pixelVec_1_0_13 = tmp_pixelVec_1_0_0_1[111 : 104];
  assign pixelVec_1_0_14 = tmp_pixelVec_1_0_0_1[119 : 112];
  assign pixelVec_1_0_15 = tmp_pixelVec_1_0_0_1[127 : 120];
  assign tmp_pixelVec_1_1_0 = tmp_pixelVec_1_0_0[255 : 128];
  assign pixelVec_1_1_0 = tmp_pixelVec_1_1_0[7 : 0];
  assign pixelVec_1_1_1 = tmp_pixelVec_1_1_0[15 : 8];
  assign pixelVec_1_1_2 = tmp_pixelVec_1_1_0[23 : 16];
  assign pixelVec_1_1_3 = tmp_pixelVec_1_1_0[31 : 24];
  assign pixelVec_1_1_4 = tmp_pixelVec_1_1_0[39 : 32];
  assign pixelVec_1_1_5 = tmp_pixelVec_1_1_0[47 : 40];
  assign pixelVec_1_1_6 = tmp_pixelVec_1_1_0[55 : 48];
  assign pixelVec_1_1_7 = tmp_pixelVec_1_1_0[63 : 56];
  assign pixelVec_1_1_8 = tmp_pixelVec_1_1_0[71 : 64];
  assign pixelVec_1_1_9 = tmp_pixelVec_1_1_0[79 : 72];
  assign pixelVec_1_1_10 = tmp_pixelVec_1_1_0[87 : 80];
  assign pixelVec_1_1_11 = tmp_pixelVec_1_1_0[95 : 88];
  assign pixelVec_1_1_12 = tmp_pixelVec_1_1_0[103 : 96];
  assign pixelVec_1_1_13 = tmp_pixelVec_1_1_0[111 : 104];
  assign pixelVec_1_1_14 = tmp_pixelVec_1_1_0[119 : 112];
  assign pixelVec_1_1_15 = tmp_pixelVec_1_1_0[127 : 120];
  assign bridge_payload_endOfPack = videoIn_payload_endOfPack;
  assign bridge_payload_frame_endOfFrame = videoIn_payload_frame_endOfFrame;
  assign bridge_payload_frame_line_endOfLine = videoIn_payload_frame_line_endOfLine;
  assign bridge_payload_frame_line_pixel_0_0_0 = pixelVec_0_0_0;
  assign bridge_payload_frame_line_pixel_0_0_1 = pixelVec_0_0_1;
  assign bridge_payload_frame_line_pixel_0_0_2 = pixelVec_0_0_2;
  assign bridge_payload_frame_line_pixel_0_0_3 = pixelVec_0_0_3;
  assign bridge_payload_frame_line_pixel_0_0_4 = pixelVec_0_0_4;
  assign bridge_payload_frame_line_pixel_0_0_5 = pixelVec_0_0_5;
  assign bridge_payload_frame_line_pixel_0_0_6 = pixelVec_0_0_6;
  assign bridge_payload_frame_line_pixel_0_0_7 = pixelVec_0_0_7;
  assign bridge_payload_frame_line_pixel_0_0_8 = pixelVec_0_0_8;
  assign bridge_payload_frame_line_pixel_0_0_9 = pixelVec_0_0_9;
  assign bridge_payload_frame_line_pixel_0_0_10 = pixelVec_0_0_10;
  assign bridge_payload_frame_line_pixel_0_0_11 = pixelVec_0_0_11;
  assign bridge_payload_frame_line_pixel_0_0_12 = pixelVec_0_0_12;
  assign bridge_payload_frame_line_pixel_0_0_13 = pixelVec_0_0_13;
  assign bridge_payload_frame_line_pixel_0_0_14 = pixelVec_0_0_14;
  assign bridge_payload_frame_line_pixel_0_0_15 = pixelVec_0_0_15;
  assign bridge_payload_frame_line_pixel_0_1_0 = pixelVec_0_1_0;
  assign bridge_payload_frame_line_pixel_0_1_1 = pixelVec_0_1_1;
  assign bridge_payload_frame_line_pixel_0_1_2 = pixelVec_0_1_2;
  assign bridge_payload_frame_line_pixel_0_1_3 = pixelVec_0_1_3;
  assign bridge_payload_frame_line_pixel_0_1_4 = pixelVec_0_1_4;
  assign bridge_payload_frame_line_pixel_0_1_5 = pixelVec_0_1_5;
  assign bridge_payload_frame_line_pixel_0_1_6 = pixelVec_0_1_6;
  assign bridge_payload_frame_line_pixel_0_1_7 = pixelVec_0_1_7;
  assign bridge_payload_frame_line_pixel_0_1_8 = pixelVec_0_1_8;
  assign bridge_payload_frame_line_pixel_0_1_9 = pixelVec_0_1_9;
  assign bridge_payload_frame_line_pixel_0_1_10 = pixelVec_0_1_10;
  assign bridge_payload_frame_line_pixel_0_1_11 = pixelVec_0_1_11;
  assign bridge_payload_frame_line_pixel_0_1_12 = pixelVec_0_1_12;
  assign bridge_payload_frame_line_pixel_0_1_13 = pixelVec_0_1_13;
  assign bridge_payload_frame_line_pixel_0_1_14 = pixelVec_0_1_14;
  assign bridge_payload_frame_line_pixel_0_1_15 = pixelVec_0_1_15;
  assign bridge_payload_frame_line_pixel_1_0_0 = pixelVec_1_0_0;
  assign bridge_payload_frame_line_pixel_1_0_1 = pixelVec_1_0_1;
  assign bridge_payload_frame_line_pixel_1_0_2 = pixelVec_1_0_2;
  assign bridge_payload_frame_line_pixel_1_0_3 = pixelVec_1_0_3;
  assign bridge_payload_frame_line_pixel_1_0_4 = pixelVec_1_0_4;
  assign bridge_payload_frame_line_pixel_1_0_5 = pixelVec_1_0_5;
  assign bridge_payload_frame_line_pixel_1_0_6 = pixelVec_1_0_6;
  assign bridge_payload_frame_line_pixel_1_0_7 = pixelVec_1_0_7;
  assign bridge_payload_frame_line_pixel_1_0_8 = pixelVec_1_0_8;
  assign bridge_payload_frame_line_pixel_1_0_9 = pixelVec_1_0_9;
  assign bridge_payload_frame_line_pixel_1_0_10 = pixelVec_1_0_10;
  assign bridge_payload_frame_line_pixel_1_0_11 = pixelVec_1_0_11;
  assign bridge_payload_frame_line_pixel_1_0_12 = pixelVec_1_0_12;
  assign bridge_payload_frame_line_pixel_1_0_13 = pixelVec_1_0_13;
  assign bridge_payload_frame_line_pixel_1_0_14 = pixelVec_1_0_14;
  assign bridge_payload_frame_line_pixel_1_0_15 = pixelVec_1_0_15;
  assign bridge_payload_frame_line_pixel_1_1_0 = pixelVec_1_1_0;
  assign bridge_payload_frame_line_pixel_1_1_1 = pixelVec_1_1_1;
  assign bridge_payload_frame_line_pixel_1_1_2 = pixelVec_1_1_2;
  assign bridge_payload_frame_line_pixel_1_1_3 = pixelVec_1_1_3;
  assign bridge_payload_frame_line_pixel_1_1_4 = pixelVec_1_1_4;
  assign bridge_payload_frame_line_pixel_1_1_5 = pixelVec_1_1_5;
  assign bridge_payload_frame_line_pixel_1_1_6 = pixelVec_1_1_6;
  assign bridge_payload_frame_line_pixel_1_1_7 = pixelVec_1_1_7;
  assign bridge_payload_frame_line_pixel_1_1_8 = pixelVec_1_1_8;
  assign bridge_payload_frame_line_pixel_1_1_9 = pixelVec_1_1_9;
  assign bridge_payload_frame_line_pixel_1_1_10 = pixelVec_1_1_10;
  assign bridge_payload_frame_line_pixel_1_1_11 = pixelVec_1_1_11;
  assign bridge_payload_frame_line_pixel_1_1_12 = pixelVec_1_1_12;
  assign bridge_payload_frame_line_pixel_1_1_13 = pixelVec_1_1_13;
  assign bridge_payload_frame_line_pixel_1_1_14 = pixelVec_1_1_14;
  assign bridge_payload_frame_line_pixel_1_1_15 = pixelVec_1_1_15;
  always @(*) begin
    bridge_thrown_valid = bridge_valid;
    if(pixelCntWontOverflowIfInc) begin
      bridge_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    bridge_ready = bridge_thrown_ready;
    if(pixelCntWontOverflowIfInc) begin
      bridge_ready = 1'b1;
    end
  end

  assign bridge_thrown_payload_frame_line_pixel_0_0_0 = bridge_payload_frame_line_pixel_0_0_0;
  assign bridge_thrown_payload_frame_line_pixel_0_0_1 = bridge_payload_frame_line_pixel_0_0_1;
  assign bridge_thrown_payload_frame_line_pixel_0_0_2 = bridge_payload_frame_line_pixel_0_0_2;
  assign bridge_thrown_payload_frame_line_pixel_0_0_3 = bridge_payload_frame_line_pixel_0_0_3;
  assign bridge_thrown_payload_frame_line_pixel_0_0_4 = bridge_payload_frame_line_pixel_0_0_4;
  assign bridge_thrown_payload_frame_line_pixel_0_0_5 = bridge_payload_frame_line_pixel_0_0_5;
  assign bridge_thrown_payload_frame_line_pixel_0_0_6 = bridge_payload_frame_line_pixel_0_0_6;
  assign bridge_thrown_payload_frame_line_pixel_0_0_7 = bridge_payload_frame_line_pixel_0_0_7;
  assign bridge_thrown_payload_frame_line_pixel_0_0_8 = bridge_payload_frame_line_pixel_0_0_8;
  assign bridge_thrown_payload_frame_line_pixel_0_0_9 = bridge_payload_frame_line_pixel_0_0_9;
  assign bridge_thrown_payload_frame_line_pixel_0_0_10 = bridge_payload_frame_line_pixel_0_0_10;
  assign bridge_thrown_payload_frame_line_pixel_0_0_11 = bridge_payload_frame_line_pixel_0_0_11;
  assign bridge_thrown_payload_frame_line_pixel_0_0_12 = bridge_payload_frame_line_pixel_0_0_12;
  assign bridge_thrown_payload_frame_line_pixel_0_0_13 = bridge_payload_frame_line_pixel_0_0_13;
  assign bridge_thrown_payload_frame_line_pixel_0_0_14 = bridge_payload_frame_line_pixel_0_0_14;
  assign bridge_thrown_payload_frame_line_pixel_0_0_15 = bridge_payload_frame_line_pixel_0_0_15;
  assign bridge_thrown_payload_frame_line_pixel_0_1_0 = bridge_payload_frame_line_pixel_0_1_0;
  assign bridge_thrown_payload_frame_line_pixel_0_1_1 = bridge_payload_frame_line_pixel_0_1_1;
  assign bridge_thrown_payload_frame_line_pixel_0_1_2 = bridge_payload_frame_line_pixel_0_1_2;
  assign bridge_thrown_payload_frame_line_pixel_0_1_3 = bridge_payload_frame_line_pixel_0_1_3;
  assign bridge_thrown_payload_frame_line_pixel_0_1_4 = bridge_payload_frame_line_pixel_0_1_4;
  assign bridge_thrown_payload_frame_line_pixel_0_1_5 = bridge_payload_frame_line_pixel_0_1_5;
  assign bridge_thrown_payload_frame_line_pixel_0_1_6 = bridge_payload_frame_line_pixel_0_1_6;
  assign bridge_thrown_payload_frame_line_pixel_0_1_7 = bridge_payload_frame_line_pixel_0_1_7;
  assign bridge_thrown_payload_frame_line_pixel_0_1_8 = bridge_payload_frame_line_pixel_0_1_8;
  assign bridge_thrown_payload_frame_line_pixel_0_1_9 = bridge_payload_frame_line_pixel_0_1_9;
  assign bridge_thrown_payload_frame_line_pixel_0_1_10 = bridge_payload_frame_line_pixel_0_1_10;
  assign bridge_thrown_payload_frame_line_pixel_0_1_11 = bridge_payload_frame_line_pixel_0_1_11;
  assign bridge_thrown_payload_frame_line_pixel_0_1_12 = bridge_payload_frame_line_pixel_0_1_12;
  assign bridge_thrown_payload_frame_line_pixel_0_1_13 = bridge_payload_frame_line_pixel_0_1_13;
  assign bridge_thrown_payload_frame_line_pixel_0_1_14 = bridge_payload_frame_line_pixel_0_1_14;
  assign bridge_thrown_payload_frame_line_pixel_0_1_15 = bridge_payload_frame_line_pixel_0_1_15;
  assign bridge_thrown_payload_frame_line_pixel_1_0_0 = bridge_payload_frame_line_pixel_1_0_0;
  assign bridge_thrown_payload_frame_line_pixel_1_0_1 = bridge_payload_frame_line_pixel_1_0_1;
  assign bridge_thrown_payload_frame_line_pixel_1_0_2 = bridge_payload_frame_line_pixel_1_0_2;
  assign bridge_thrown_payload_frame_line_pixel_1_0_3 = bridge_payload_frame_line_pixel_1_0_3;
  assign bridge_thrown_payload_frame_line_pixel_1_0_4 = bridge_payload_frame_line_pixel_1_0_4;
  assign bridge_thrown_payload_frame_line_pixel_1_0_5 = bridge_payload_frame_line_pixel_1_0_5;
  assign bridge_thrown_payload_frame_line_pixel_1_0_6 = bridge_payload_frame_line_pixel_1_0_6;
  assign bridge_thrown_payload_frame_line_pixel_1_0_7 = bridge_payload_frame_line_pixel_1_0_7;
  assign bridge_thrown_payload_frame_line_pixel_1_0_8 = bridge_payload_frame_line_pixel_1_0_8;
  assign bridge_thrown_payload_frame_line_pixel_1_0_9 = bridge_payload_frame_line_pixel_1_0_9;
  assign bridge_thrown_payload_frame_line_pixel_1_0_10 = bridge_payload_frame_line_pixel_1_0_10;
  assign bridge_thrown_payload_frame_line_pixel_1_0_11 = bridge_payload_frame_line_pixel_1_0_11;
  assign bridge_thrown_payload_frame_line_pixel_1_0_12 = bridge_payload_frame_line_pixel_1_0_12;
  assign bridge_thrown_payload_frame_line_pixel_1_0_13 = bridge_payload_frame_line_pixel_1_0_13;
  assign bridge_thrown_payload_frame_line_pixel_1_0_14 = bridge_payload_frame_line_pixel_1_0_14;
  assign bridge_thrown_payload_frame_line_pixel_1_0_15 = bridge_payload_frame_line_pixel_1_0_15;
  assign bridge_thrown_payload_frame_line_pixel_1_1_0 = bridge_payload_frame_line_pixel_1_1_0;
  assign bridge_thrown_payload_frame_line_pixel_1_1_1 = bridge_payload_frame_line_pixel_1_1_1;
  assign bridge_thrown_payload_frame_line_pixel_1_1_2 = bridge_payload_frame_line_pixel_1_1_2;
  assign bridge_thrown_payload_frame_line_pixel_1_1_3 = bridge_payload_frame_line_pixel_1_1_3;
  assign bridge_thrown_payload_frame_line_pixel_1_1_4 = bridge_payload_frame_line_pixel_1_1_4;
  assign bridge_thrown_payload_frame_line_pixel_1_1_5 = bridge_payload_frame_line_pixel_1_1_5;
  assign bridge_thrown_payload_frame_line_pixel_1_1_6 = bridge_payload_frame_line_pixel_1_1_6;
  assign bridge_thrown_payload_frame_line_pixel_1_1_7 = bridge_payload_frame_line_pixel_1_1_7;
  assign bridge_thrown_payload_frame_line_pixel_1_1_8 = bridge_payload_frame_line_pixel_1_1_8;
  assign bridge_thrown_payload_frame_line_pixel_1_1_9 = bridge_payload_frame_line_pixel_1_1_9;
  assign bridge_thrown_payload_frame_line_pixel_1_1_10 = bridge_payload_frame_line_pixel_1_1_10;
  assign bridge_thrown_payload_frame_line_pixel_1_1_11 = bridge_payload_frame_line_pixel_1_1_11;
  assign bridge_thrown_payload_frame_line_pixel_1_1_12 = bridge_payload_frame_line_pixel_1_1_12;
  assign bridge_thrown_payload_frame_line_pixel_1_1_13 = bridge_payload_frame_line_pixel_1_1_13;
  assign bridge_thrown_payload_frame_line_pixel_1_1_14 = bridge_payload_frame_line_pixel_1_1_14;
  assign bridge_thrown_payload_frame_line_pixel_1_1_15 = bridge_payload_frame_line_pixel_1_1_15;
  assign bridge_thrown_payload_frame_line_endOfLine = bridge_payload_frame_line_endOfLine;
  assign bridge_thrown_payload_frame_endOfFrame = bridge_payload_frame_endOfFrame;
  assign bridge_thrown_payload_endOfPack = bridge_payload_endOfPack;
  assign videoOut_valid = bridge_thrown_valid;
  assign bridge_thrown_ready = videoOut_ready;
  assign videoOut_payload_frame_line_pixel_0_0_0 = bridge_thrown_payload_frame_line_pixel_0_0_0;
  assign videoOut_payload_frame_line_pixel_0_0_1 = bridge_thrown_payload_frame_line_pixel_0_0_1;
  assign videoOut_payload_frame_line_pixel_0_0_2 = bridge_thrown_payload_frame_line_pixel_0_0_2;
  assign videoOut_payload_frame_line_pixel_0_0_3 = bridge_thrown_payload_frame_line_pixel_0_0_3;
  assign videoOut_payload_frame_line_pixel_0_0_4 = bridge_thrown_payload_frame_line_pixel_0_0_4;
  assign videoOut_payload_frame_line_pixel_0_0_5 = bridge_thrown_payload_frame_line_pixel_0_0_5;
  assign videoOut_payload_frame_line_pixel_0_0_6 = bridge_thrown_payload_frame_line_pixel_0_0_6;
  assign videoOut_payload_frame_line_pixel_0_0_7 = bridge_thrown_payload_frame_line_pixel_0_0_7;
  assign videoOut_payload_frame_line_pixel_0_0_8 = bridge_thrown_payload_frame_line_pixel_0_0_8;
  assign videoOut_payload_frame_line_pixel_0_0_9 = bridge_thrown_payload_frame_line_pixel_0_0_9;
  assign videoOut_payload_frame_line_pixel_0_0_10 = bridge_thrown_payload_frame_line_pixel_0_0_10;
  assign videoOut_payload_frame_line_pixel_0_0_11 = bridge_thrown_payload_frame_line_pixel_0_0_11;
  assign videoOut_payload_frame_line_pixel_0_0_12 = bridge_thrown_payload_frame_line_pixel_0_0_12;
  assign videoOut_payload_frame_line_pixel_0_0_13 = bridge_thrown_payload_frame_line_pixel_0_0_13;
  assign videoOut_payload_frame_line_pixel_0_0_14 = bridge_thrown_payload_frame_line_pixel_0_0_14;
  assign videoOut_payload_frame_line_pixel_0_0_15 = bridge_thrown_payload_frame_line_pixel_0_0_15;
  assign videoOut_payload_frame_line_pixel_0_1_0 = bridge_thrown_payload_frame_line_pixel_0_1_0;
  assign videoOut_payload_frame_line_pixel_0_1_1 = bridge_thrown_payload_frame_line_pixel_0_1_1;
  assign videoOut_payload_frame_line_pixel_0_1_2 = bridge_thrown_payload_frame_line_pixel_0_1_2;
  assign videoOut_payload_frame_line_pixel_0_1_3 = bridge_thrown_payload_frame_line_pixel_0_1_3;
  assign videoOut_payload_frame_line_pixel_0_1_4 = bridge_thrown_payload_frame_line_pixel_0_1_4;
  assign videoOut_payload_frame_line_pixel_0_1_5 = bridge_thrown_payload_frame_line_pixel_0_1_5;
  assign videoOut_payload_frame_line_pixel_0_1_6 = bridge_thrown_payload_frame_line_pixel_0_1_6;
  assign videoOut_payload_frame_line_pixel_0_1_7 = bridge_thrown_payload_frame_line_pixel_0_1_7;
  assign videoOut_payload_frame_line_pixel_0_1_8 = bridge_thrown_payload_frame_line_pixel_0_1_8;
  assign videoOut_payload_frame_line_pixel_0_1_9 = bridge_thrown_payload_frame_line_pixel_0_1_9;
  assign videoOut_payload_frame_line_pixel_0_1_10 = bridge_thrown_payload_frame_line_pixel_0_1_10;
  assign videoOut_payload_frame_line_pixel_0_1_11 = bridge_thrown_payload_frame_line_pixel_0_1_11;
  assign videoOut_payload_frame_line_pixel_0_1_12 = bridge_thrown_payload_frame_line_pixel_0_1_12;
  assign videoOut_payload_frame_line_pixel_0_1_13 = bridge_thrown_payload_frame_line_pixel_0_1_13;
  assign videoOut_payload_frame_line_pixel_0_1_14 = bridge_thrown_payload_frame_line_pixel_0_1_14;
  assign videoOut_payload_frame_line_pixel_0_1_15 = bridge_thrown_payload_frame_line_pixel_0_1_15;
  assign videoOut_payload_frame_line_pixel_1_0_0 = bridge_thrown_payload_frame_line_pixel_1_0_0;
  assign videoOut_payload_frame_line_pixel_1_0_1 = bridge_thrown_payload_frame_line_pixel_1_0_1;
  assign videoOut_payload_frame_line_pixel_1_0_2 = bridge_thrown_payload_frame_line_pixel_1_0_2;
  assign videoOut_payload_frame_line_pixel_1_0_3 = bridge_thrown_payload_frame_line_pixel_1_0_3;
  assign videoOut_payload_frame_line_pixel_1_0_4 = bridge_thrown_payload_frame_line_pixel_1_0_4;
  assign videoOut_payload_frame_line_pixel_1_0_5 = bridge_thrown_payload_frame_line_pixel_1_0_5;
  assign videoOut_payload_frame_line_pixel_1_0_6 = bridge_thrown_payload_frame_line_pixel_1_0_6;
  assign videoOut_payload_frame_line_pixel_1_0_7 = bridge_thrown_payload_frame_line_pixel_1_0_7;
  assign videoOut_payload_frame_line_pixel_1_0_8 = bridge_thrown_payload_frame_line_pixel_1_0_8;
  assign videoOut_payload_frame_line_pixel_1_0_9 = bridge_thrown_payload_frame_line_pixel_1_0_9;
  assign videoOut_payload_frame_line_pixel_1_0_10 = bridge_thrown_payload_frame_line_pixel_1_0_10;
  assign videoOut_payload_frame_line_pixel_1_0_11 = bridge_thrown_payload_frame_line_pixel_1_0_11;
  assign videoOut_payload_frame_line_pixel_1_0_12 = bridge_thrown_payload_frame_line_pixel_1_0_12;
  assign videoOut_payload_frame_line_pixel_1_0_13 = bridge_thrown_payload_frame_line_pixel_1_0_13;
  assign videoOut_payload_frame_line_pixel_1_0_14 = bridge_thrown_payload_frame_line_pixel_1_0_14;
  assign videoOut_payload_frame_line_pixel_1_0_15 = bridge_thrown_payload_frame_line_pixel_1_0_15;
  assign videoOut_payload_frame_line_pixel_1_1_0 = bridge_thrown_payload_frame_line_pixel_1_1_0;
  assign videoOut_payload_frame_line_pixel_1_1_1 = bridge_thrown_payload_frame_line_pixel_1_1_1;
  assign videoOut_payload_frame_line_pixel_1_1_2 = bridge_thrown_payload_frame_line_pixel_1_1_2;
  assign videoOut_payload_frame_line_pixel_1_1_3 = bridge_thrown_payload_frame_line_pixel_1_1_3;
  assign videoOut_payload_frame_line_pixel_1_1_4 = bridge_thrown_payload_frame_line_pixel_1_1_4;
  assign videoOut_payload_frame_line_pixel_1_1_5 = bridge_thrown_payload_frame_line_pixel_1_1_5;
  assign videoOut_payload_frame_line_pixel_1_1_6 = bridge_thrown_payload_frame_line_pixel_1_1_6;
  assign videoOut_payload_frame_line_pixel_1_1_7 = bridge_thrown_payload_frame_line_pixel_1_1_7;
  assign videoOut_payload_frame_line_pixel_1_1_8 = bridge_thrown_payload_frame_line_pixel_1_1_8;
  assign videoOut_payload_frame_line_pixel_1_1_9 = bridge_thrown_payload_frame_line_pixel_1_1_9;
  assign videoOut_payload_frame_line_pixel_1_1_10 = bridge_thrown_payload_frame_line_pixel_1_1_10;
  assign videoOut_payload_frame_line_pixel_1_1_11 = bridge_thrown_payload_frame_line_pixel_1_1_11;
  assign videoOut_payload_frame_line_pixel_1_1_12 = bridge_thrown_payload_frame_line_pixel_1_1_12;
  assign videoOut_payload_frame_line_pixel_1_1_13 = bridge_thrown_payload_frame_line_pixel_1_1_13;
  assign videoOut_payload_frame_line_pixel_1_1_14 = bridge_thrown_payload_frame_line_pixel_1_1_14;
  assign videoOut_payload_frame_line_pixel_1_1_15 = bridge_thrown_payload_frame_line_pixel_1_1_15;
  assign videoOut_payload_frame_line_endOfLine = bridge_thrown_payload_frame_line_endOfLine;
  assign videoOut_payload_frame_endOfFrame = bridge_thrown_payload_frame_endOfFrame;
  assign videoOut_payload_endOfPack = bridge_thrown_payload_endOfPack;
  always @(posedge clk) begin
    if(videoInFire) begin
      pixelBuffer <= {{videoIn_payload_frame_line_pixel_1_15,{videoIn_payload_frame_line_pixel_1_14,{videoIn_payload_frame_line_pixel_1_13,{videoIn_payload_frame_line_pixel_1_12,{videoIn_payload_frame_line_pixel_1_11,{videoIn_payload_frame_line_pixel_1_10,{videoIn_payload_frame_line_pixel_1_9,{tmp_pixelBuffer,tmp_pixelBuffer_1}}}}}}}},{videoIn_payload_frame_line_pixel_0_15,{videoIn_payload_frame_line_pixel_0_14,{videoIn_payload_frame_line_pixel_0_13,{videoIn_payload_frame_line_pixel_0_12,{videoIn_payload_frame_line_pixel_0_11,{videoIn_payload_frame_line_pixel_0_10,{videoIn_payload_frame_line_pixel_0_9,{tmp_pixelBuffer_2,tmp_pixelBuffer_3}}}}}}}}};
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      pixelCnt_value <= 1'b0;
    end else begin
      pixelCnt_value <= pixelCnt_valueNext;
    end
  end


endmodule

module LineBufferValid (
  input               videoIn_valid,
  output              videoIn_ready,
  input      [7:0]    videoIn_payload_frame_line_pixel_0,
  input      [7:0]    videoIn_payload_frame_line_pixel_1,
  input      [7:0]    videoIn_payload_frame_line_pixel_2,
  input      [7:0]    videoIn_payload_frame_line_pixel_3,
  input      [7:0]    videoIn_payload_frame_line_pixel_4,
  input      [7:0]    videoIn_payload_frame_line_pixel_5,
  input      [7:0]    videoIn_payload_frame_line_pixel_6,
  input      [7:0]    videoIn_payload_frame_line_pixel_7,
  input      [7:0]    videoIn_payload_frame_line_pixel_8,
  input      [7:0]    videoIn_payload_frame_line_pixel_9,
  input      [7:0]    videoIn_payload_frame_line_pixel_10,
  input      [7:0]    videoIn_payload_frame_line_pixel_11,
  input      [7:0]    videoIn_payload_frame_line_pixel_12,
  input      [7:0]    videoIn_payload_frame_line_pixel_13,
  input      [7:0]    videoIn_payload_frame_line_pixel_14,
  input      [7:0]    videoIn_payload_frame_line_pixel_15,
  input               videoIn_payload_frame_line_endOfLine,
  input               videoIn_payload_frame_endOfFrame,
  input               videoIn_payload_endOfPack,
  output              videoOut_valid,
  input               videoOut_ready,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_0_15,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_0,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_1,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_2,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_3,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_4,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_5,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_6,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_7,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_8,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_9,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_10,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_11,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_12,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_13,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_14,
  output     [7:0]    videoOut_payload_frame_line_pixel_1_15,
  output              videoOut_payload_frame_line_endOfLine,
  output              videoOut_payload_frame_endOfFrame,
  output              videoOut_payload_endOfPack,
  input               clk,
  input               reset
);

  wire                fifo_flush;
  reg                 videoIn_fork_io_outputs_1_ready;
  reg                 fifo_pop_fork_io_outputs_0_ready;
  wire                fifo_push_ready;
  wire                fifo_pop_valid;
  wire       [7:0]    fifo_pop_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_payload_0_pixel_15;
  wire                fifo_pop_payload_0_endOfLine;
  wire                videoIn_fork_io_input_ready;
  wire                videoIn_fork_io_outputs_0_valid;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_0;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_1;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_2;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_3;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_4;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_5;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_6;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_7;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_8;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_9;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_10;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_11;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_12;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_13;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_14;
  wire       [7:0]    videoIn_fork_io_outputs_0_payload_frame_line_pixel_15;
  wire                videoIn_fork_io_outputs_0_payload_frame_line_endOfLine;
  wire                videoIn_fork_io_outputs_0_payload_frame_endOfFrame;
  wire                videoIn_fork_io_outputs_0_payload_endOfPack;
  wire                videoIn_fork_io_outputs_1_valid;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_0;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_1;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_2;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_3;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_4;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_5;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_6;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_7;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_8;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_9;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_10;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_11;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_12;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_13;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_14;
  wire       [7:0]    videoIn_fork_io_outputs_1_payload_frame_line_pixel_15;
  wire                videoIn_fork_io_outputs_1_payload_frame_line_endOfLine;
  wire                videoIn_fork_io_outputs_1_payload_frame_endOfFrame;
  wire                videoIn_fork_io_outputs_1_payload_endOfPack;
  wire                fifo_pop_fork_io_input_ready;
  wire                fifo_pop_fork_io_outputs_0_valid;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_0_payload_0_pixel_15;
  wire                fifo_pop_fork_io_outputs_0_payload_0_endOfLine;
  wire                fifo_pop_fork_io_outputs_1_valid;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_0;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_1;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_2;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_3;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_4;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_5;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_6;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_7;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_8;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_9;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_10;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_11;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_12;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_13;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_14;
  wire       [7:0]    fifo_pop_fork_io_outputs_1_payload_0_pixel_15;
  wire                fifo_pop_fork_io_outputs_1_payload_0_endOfLine;
  wire                in2outThrowCond;
  wire                feedbackAddCond;
  reg                 in2outThrown_valid;
  wire                in2outThrown_ready;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_0;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_1;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_2;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_3;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_4;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_5;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_6;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_7;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_8;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_9;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_10;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_11;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_12;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_13;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_14;
  wire       [7:0]    in2outThrown_payload_frame_line_pixel_15;
  wire                in2outThrown_payload_frame_line_endOfLine;
  wire                in2outThrown_payload_frame_endOfFrame;
  wire                in2outThrown_payload_endOfPack;
  reg                 feedbackAdded_valid;
  wire                feedbackAdded_ready;
  wire       [7:0]    feedbackAdded_payload_0_pixel_0;
  wire       [7:0]    feedbackAdded_payload_0_pixel_1;
  wire       [7:0]    feedbackAdded_payload_0_pixel_2;
  wire       [7:0]    feedbackAdded_payload_0_pixel_3;
  wire       [7:0]    feedbackAdded_payload_0_pixel_4;
  wire       [7:0]    feedbackAdded_payload_0_pixel_5;
  wire       [7:0]    feedbackAdded_payload_0_pixel_6;
  wire       [7:0]    feedbackAdded_payload_0_pixel_7;
  wire       [7:0]    feedbackAdded_payload_0_pixel_8;
  wire       [7:0]    feedbackAdded_payload_0_pixel_9;
  wire       [7:0]    feedbackAdded_payload_0_pixel_10;
  wire       [7:0]    feedbackAdded_payload_0_pixel_11;
  wire       [7:0]    feedbackAdded_payload_0_pixel_12;
  wire       [7:0]    feedbackAdded_payload_0_pixel_13;
  wire       [7:0]    feedbackAdded_payload_0_pixel_14;
  wire       [7:0]    feedbackAdded_payload_0_pixel_15;
  wire                feedbackAdded_payload_0_endOfLine;
  wire                in2fifoJoinFeedback_valid;
  wire                in2fifoJoinFeedback_ready;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_0;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_1;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_2;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_3;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_4;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_5;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_6;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_7;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_8;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_9;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_10;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_11;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_12;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_13;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_14;
  wire       [7:0]    in2fifoJoinFeedback_payload__1_frame_line_pixel_15;
  wire                in2fifoJoinFeedback_payload__1_frame_line_endOfLine;
  wire                in2fifoJoinFeedback_payload__1_frame_endOfFrame;
  wire                in2fifoJoinFeedback_payload__1_endOfPack;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_0;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_1;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_2;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_3;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_4;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_5;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_6;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_7;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_8;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_9;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_10;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_11;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_12;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_13;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_14;
  wire       [7:0]    in2fifoJoinFeedback_payload__2_0_pixel_15;
  wire                in2fifoJoinFeedback_payload__2_0_endOfLine;
  wire                in2fifoJoinFeedback_fire;
  wire                in2fifoJoinFeedback_fire_1;
  wire                in2outJoinFifo2out_valid;
  wire                in2outJoinFifo2out_ready;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_0;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_1;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_2;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_3;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_4;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_5;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_6;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_7;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_8;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_9;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_10;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_11;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_12;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_13;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_14;
  wire       [7:0]    in2outJoinFifo2out_payload__1_frame_line_pixel_15;
  wire                in2outJoinFifo2out_payload__1_frame_line_endOfLine;
  wire                in2outJoinFifo2out_payload__1_frame_endOfFrame;
  wire                in2outJoinFifo2out_payload__1_endOfPack;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_0;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_1;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_2;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_3;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_4;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_5;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_6;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_7;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_8;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_9;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_10;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_11;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_12;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_13;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_14;
  wire       [7:0]    in2outJoinFifo2out_payload__2_0_pixel_15;
  wire                in2outJoinFifo2out_payload__2_0_endOfLine;
  wire                in2outJoinFifo2out_fire;
  wire                in2outJoinFifo2out_fire_1;
  wire                ioVideoInFire;
  reg                 lineCnt_willIncrement;
  reg                 lineCnt_willClear;
  reg        [0:0]    lineCnt_valueNext;
  reg        [0:0]    lineCnt_value;
  wire                lineCnt_willOverflowIfInc;
  wire                lineCnt_willOverflow;
  wire                lineCntWontOverflowIfInc;
  wire                when_LineBufferValid_l58;
  wire                when_LineBufferValid_l59;

  StreamFifoHighPerf fifo (
    .push_valid                  (in2fifoJoinFeedback_valid                                ), //i
    .push_ready                  (fifo_push_ready                                          ), //o
    .push_payload_0_pixel_0      (in2fifoJoinFeedback_payload__1_frame_line_pixel_0[7:0]   ), //i
    .push_payload_0_pixel_1      (in2fifoJoinFeedback_payload__1_frame_line_pixel_1[7:0]   ), //i
    .push_payload_0_pixel_2      (in2fifoJoinFeedback_payload__1_frame_line_pixel_2[7:0]   ), //i
    .push_payload_0_pixel_3      (in2fifoJoinFeedback_payload__1_frame_line_pixel_3[7:0]   ), //i
    .push_payload_0_pixel_4      (in2fifoJoinFeedback_payload__1_frame_line_pixel_4[7:0]   ), //i
    .push_payload_0_pixel_5      (in2fifoJoinFeedback_payload__1_frame_line_pixel_5[7:0]   ), //i
    .push_payload_0_pixel_6      (in2fifoJoinFeedback_payload__1_frame_line_pixel_6[7:0]   ), //i
    .push_payload_0_pixel_7      (in2fifoJoinFeedback_payload__1_frame_line_pixel_7[7:0]   ), //i
    .push_payload_0_pixel_8      (in2fifoJoinFeedback_payload__1_frame_line_pixel_8[7:0]   ), //i
    .push_payload_0_pixel_9      (in2fifoJoinFeedback_payload__1_frame_line_pixel_9[7:0]   ), //i
    .push_payload_0_pixel_10     (in2fifoJoinFeedback_payload__1_frame_line_pixel_10[7:0]  ), //i
    .push_payload_0_pixel_11     (in2fifoJoinFeedback_payload__1_frame_line_pixel_11[7:0]  ), //i
    .push_payload_0_pixel_12     (in2fifoJoinFeedback_payload__1_frame_line_pixel_12[7:0]  ), //i
    .push_payload_0_pixel_13     (in2fifoJoinFeedback_payload__1_frame_line_pixel_13[7:0]  ), //i
    .push_payload_0_pixel_14     (in2fifoJoinFeedback_payload__1_frame_line_pixel_14[7:0]  ), //i
    .push_payload_0_pixel_15     (in2fifoJoinFeedback_payload__1_frame_line_pixel_15[7:0]  ), //i
    .push_payload_0_endOfLine    (in2fifoJoinFeedback_payload__1_frame_line_endOfLine      ), //i
    .pop_valid                   (fifo_pop_valid                                           ), //o
    .pop_ready                   (fifo_pop_fork_io_input_ready                             ), //i
    .pop_payload_0_pixel_0       (fifo_pop_payload_0_pixel_0[7:0]                          ), //o
    .pop_payload_0_pixel_1       (fifo_pop_payload_0_pixel_1[7:0]                          ), //o
    .pop_payload_0_pixel_2       (fifo_pop_payload_0_pixel_2[7:0]                          ), //o
    .pop_payload_0_pixel_3       (fifo_pop_payload_0_pixel_3[7:0]                          ), //o
    .pop_payload_0_pixel_4       (fifo_pop_payload_0_pixel_4[7:0]                          ), //o
    .pop_payload_0_pixel_5       (fifo_pop_payload_0_pixel_5[7:0]                          ), //o
    .pop_payload_0_pixel_6       (fifo_pop_payload_0_pixel_6[7:0]                          ), //o
    .pop_payload_0_pixel_7       (fifo_pop_payload_0_pixel_7[7:0]                          ), //o
    .pop_payload_0_pixel_8       (fifo_pop_payload_0_pixel_8[7:0]                          ), //o
    .pop_payload_0_pixel_9       (fifo_pop_payload_0_pixel_9[7:0]                          ), //o
    .pop_payload_0_pixel_10      (fifo_pop_payload_0_pixel_10[7:0]                         ), //o
    .pop_payload_0_pixel_11      (fifo_pop_payload_0_pixel_11[7:0]                         ), //o
    .pop_payload_0_pixel_12      (fifo_pop_payload_0_pixel_12[7:0]                         ), //o
    .pop_payload_0_pixel_13      (fifo_pop_payload_0_pixel_13[7:0]                         ), //o
    .pop_payload_0_pixel_14      (fifo_pop_payload_0_pixel_14[7:0]                         ), //o
    .pop_payload_0_pixel_15      (fifo_pop_payload_0_pixel_15[7:0]                         ), //o
    .pop_payload_0_endOfLine     (fifo_pop_payload_0_endOfLine                             ), //o
    .flush                       (fifo_flush                                               ), //i
    .clk                         (clk                                                      ), //i
    .reset                       (reset                                                    )  //i
  );
  StreamFork videoIn_fork (
    .io_input_valid                               (videoIn_valid                                               ), //i
    .io_input_ready                               (videoIn_fork_io_input_ready                                 ), //o
    .io_input_payload_frame_line_pixel_0          (videoIn_payload_frame_line_pixel_0[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_1          (videoIn_payload_frame_line_pixel_1[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_2          (videoIn_payload_frame_line_pixel_2[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_3          (videoIn_payload_frame_line_pixel_3[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_4          (videoIn_payload_frame_line_pixel_4[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_5          (videoIn_payload_frame_line_pixel_5[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_6          (videoIn_payload_frame_line_pixel_6[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_7          (videoIn_payload_frame_line_pixel_7[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_8          (videoIn_payload_frame_line_pixel_8[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_9          (videoIn_payload_frame_line_pixel_9[7:0]                     ), //i
    .io_input_payload_frame_line_pixel_10         (videoIn_payload_frame_line_pixel_10[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_11         (videoIn_payload_frame_line_pixel_11[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_12         (videoIn_payload_frame_line_pixel_12[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_13         (videoIn_payload_frame_line_pixel_13[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_14         (videoIn_payload_frame_line_pixel_14[7:0]                    ), //i
    .io_input_payload_frame_line_pixel_15         (videoIn_payload_frame_line_pixel_15[7:0]                    ), //i
    .io_input_payload_frame_line_endOfLine        (videoIn_payload_frame_line_endOfLine                        ), //i
    .io_input_payload_frame_endOfFrame            (videoIn_payload_frame_endOfFrame                            ), //i
    .io_input_payload_endOfPack                   (videoIn_payload_endOfPack                                   ), //i
    .io_outputs_0_valid                           (videoIn_fork_io_outputs_0_valid                             ), //o
    .io_outputs_0_ready                           (in2fifoJoinFeedback_fire                                    ), //i
    .io_outputs_0_payload_frame_line_pixel_0      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_1      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_2      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_3      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_4      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_5      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_6      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_7      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_8      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_9      (videoIn_fork_io_outputs_0_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_frame_line_pixel_10     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_11     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_12     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_13     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_14     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_frame_line_pixel_15     (videoIn_fork_io_outputs_0_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_frame_line_endOfLine    (videoIn_fork_io_outputs_0_payload_frame_line_endOfLine      ), //o
    .io_outputs_0_payload_frame_endOfFrame        (videoIn_fork_io_outputs_0_payload_frame_endOfFrame          ), //o
    .io_outputs_0_payload_endOfPack               (videoIn_fork_io_outputs_0_payload_endOfPack                 ), //o
    .io_outputs_1_valid                           (videoIn_fork_io_outputs_1_valid                             ), //o
    .io_outputs_1_ready                           (videoIn_fork_io_outputs_1_ready                             ), //i
    .io_outputs_1_payload_frame_line_pixel_0      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_1      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_2      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_3      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_4      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_5      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_6      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_7      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_8      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_9      (videoIn_fork_io_outputs_1_payload_frame_line_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_frame_line_pixel_10     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_11     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_12     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_13     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_14     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_frame_line_pixel_15     (videoIn_fork_io_outputs_1_payload_frame_line_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_frame_line_endOfLine    (videoIn_fork_io_outputs_1_payload_frame_line_endOfLine      ), //o
    .io_outputs_1_payload_frame_endOfFrame        (videoIn_fork_io_outputs_1_payload_frame_endOfFrame          ), //o
    .io_outputs_1_payload_endOfPack               (videoIn_fork_io_outputs_1_payload_endOfPack                 ), //o
    .clk                                          (clk                                                         ), //i
    .reset                                        (reset                                                       )  //i
  );
  StreamFork_1 fifo_pop_fork (
    .io_input_valid                      (fifo_pop_valid                                      ), //i
    .io_input_ready                      (fifo_pop_fork_io_input_ready                        ), //o
    .io_input_payload_0_pixel_0          (fifo_pop_payload_0_pixel_0[7:0]                     ), //i
    .io_input_payload_0_pixel_1          (fifo_pop_payload_0_pixel_1[7:0]                     ), //i
    .io_input_payload_0_pixel_2          (fifo_pop_payload_0_pixel_2[7:0]                     ), //i
    .io_input_payload_0_pixel_3          (fifo_pop_payload_0_pixel_3[7:0]                     ), //i
    .io_input_payload_0_pixel_4          (fifo_pop_payload_0_pixel_4[7:0]                     ), //i
    .io_input_payload_0_pixel_5          (fifo_pop_payload_0_pixel_5[7:0]                     ), //i
    .io_input_payload_0_pixel_6          (fifo_pop_payload_0_pixel_6[7:0]                     ), //i
    .io_input_payload_0_pixel_7          (fifo_pop_payload_0_pixel_7[7:0]                     ), //i
    .io_input_payload_0_pixel_8          (fifo_pop_payload_0_pixel_8[7:0]                     ), //i
    .io_input_payload_0_pixel_9          (fifo_pop_payload_0_pixel_9[7:0]                     ), //i
    .io_input_payload_0_pixel_10         (fifo_pop_payload_0_pixel_10[7:0]                    ), //i
    .io_input_payload_0_pixel_11         (fifo_pop_payload_0_pixel_11[7:0]                    ), //i
    .io_input_payload_0_pixel_12         (fifo_pop_payload_0_pixel_12[7:0]                    ), //i
    .io_input_payload_0_pixel_13         (fifo_pop_payload_0_pixel_13[7:0]                    ), //i
    .io_input_payload_0_pixel_14         (fifo_pop_payload_0_pixel_14[7:0]                    ), //i
    .io_input_payload_0_pixel_15         (fifo_pop_payload_0_pixel_15[7:0]                    ), //i
    .io_input_payload_0_endOfLine        (fifo_pop_payload_0_endOfLine                        ), //i
    .io_outputs_0_valid                  (fifo_pop_fork_io_outputs_0_valid                    ), //o
    .io_outputs_0_ready                  (fifo_pop_fork_io_outputs_0_ready                    ), //i
    .io_outputs_0_payload_0_pixel_0      (fifo_pop_fork_io_outputs_0_payload_0_pixel_0[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_1      (fifo_pop_fork_io_outputs_0_payload_0_pixel_1[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_2      (fifo_pop_fork_io_outputs_0_payload_0_pixel_2[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_3      (fifo_pop_fork_io_outputs_0_payload_0_pixel_3[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_4      (fifo_pop_fork_io_outputs_0_payload_0_pixel_4[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_5      (fifo_pop_fork_io_outputs_0_payload_0_pixel_5[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_6      (fifo_pop_fork_io_outputs_0_payload_0_pixel_6[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_7      (fifo_pop_fork_io_outputs_0_payload_0_pixel_7[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_8      (fifo_pop_fork_io_outputs_0_payload_0_pixel_8[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_9      (fifo_pop_fork_io_outputs_0_payload_0_pixel_9[7:0]   ), //o
    .io_outputs_0_payload_0_pixel_10     (fifo_pop_fork_io_outputs_0_payload_0_pixel_10[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_11     (fifo_pop_fork_io_outputs_0_payload_0_pixel_11[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_12     (fifo_pop_fork_io_outputs_0_payload_0_pixel_12[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_13     (fifo_pop_fork_io_outputs_0_payload_0_pixel_13[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_14     (fifo_pop_fork_io_outputs_0_payload_0_pixel_14[7:0]  ), //o
    .io_outputs_0_payload_0_pixel_15     (fifo_pop_fork_io_outputs_0_payload_0_pixel_15[7:0]  ), //o
    .io_outputs_0_payload_0_endOfLine    (fifo_pop_fork_io_outputs_0_payload_0_endOfLine      ), //o
    .io_outputs_1_valid                  (fifo_pop_fork_io_outputs_1_valid                    ), //o
    .io_outputs_1_ready                  (in2outJoinFifo2out_fire_1                           ), //i
    .io_outputs_1_payload_0_pixel_0      (fifo_pop_fork_io_outputs_1_payload_0_pixel_0[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_1      (fifo_pop_fork_io_outputs_1_payload_0_pixel_1[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_2      (fifo_pop_fork_io_outputs_1_payload_0_pixel_2[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_3      (fifo_pop_fork_io_outputs_1_payload_0_pixel_3[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_4      (fifo_pop_fork_io_outputs_1_payload_0_pixel_4[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_5      (fifo_pop_fork_io_outputs_1_payload_0_pixel_5[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_6      (fifo_pop_fork_io_outputs_1_payload_0_pixel_6[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_7      (fifo_pop_fork_io_outputs_1_payload_0_pixel_7[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_8      (fifo_pop_fork_io_outputs_1_payload_0_pixel_8[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_9      (fifo_pop_fork_io_outputs_1_payload_0_pixel_9[7:0]   ), //o
    .io_outputs_1_payload_0_pixel_10     (fifo_pop_fork_io_outputs_1_payload_0_pixel_10[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_11     (fifo_pop_fork_io_outputs_1_payload_0_pixel_11[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_12     (fifo_pop_fork_io_outputs_1_payload_0_pixel_12[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_13     (fifo_pop_fork_io_outputs_1_payload_0_pixel_13[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_14     (fifo_pop_fork_io_outputs_1_payload_0_pixel_14[7:0]  ), //o
    .io_outputs_1_payload_0_pixel_15     (fifo_pop_fork_io_outputs_1_payload_0_pixel_15[7:0]  ), //o
    .io_outputs_1_payload_0_endOfLine    (fifo_pop_fork_io_outputs_1_payload_0_endOfLine      ), //o
    .clk                                 (clk                                                 ), //i
    .reset                               (reset                                               )  //i
  );
  assign videoIn_ready = videoIn_fork_io_input_ready;
  always @(*) begin
    in2outThrown_valid = videoIn_fork_io_outputs_1_valid;
    if(in2outThrowCond) begin
      in2outThrown_valid = 1'b0;
    end
  end

  always @(*) begin
    videoIn_fork_io_outputs_1_ready = in2outThrown_ready;
    if(in2outThrowCond) begin
      videoIn_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign in2outThrown_payload_frame_line_pixel_0 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_0;
  assign in2outThrown_payload_frame_line_pixel_1 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_1;
  assign in2outThrown_payload_frame_line_pixel_2 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_2;
  assign in2outThrown_payload_frame_line_pixel_3 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_3;
  assign in2outThrown_payload_frame_line_pixel_4 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_4;
  assign in2outThrown_payload_frame_line_pixel_5 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_5;
  assign in2outThrown_payload_frame_line_pixel_6 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_6;
  assign in2outThrown_payload_frame_line_pixel_7 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_7;
  assign in2outThrown_payload_frame_line_pixel_8 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_8;
  assign in2outThrown_payload_frame_line_pixel_9 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_9;
  assign in2outThrown_payload_frame_line_pixel_10 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_10;
  assign in2outThrown_payload_frame_line_pixel_11 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_11;
  assign in2outThrown_payload_frame_line_pixel_12 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_12;
  assign in2outThrown_payload_frame_line_pixel_13 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_13;
  assign in2outThrown_payload_frame_line_pixel_14 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_14;
  assign in2outThrown_payload_frame_line_pixel_15 = videoIn_fork_io_outputs_1_payload_frame_line_pixel_15;
  assign in2outThrown_payload_frame_line_endOfLine = videoIn_fork_io_outputs_1_payload_frame_line_endOfLine;
  assign in2outThrown_payload_frame_endOfFrame = videoIn_fork_io_outputs_1_payload_frame_endOfFrame;
  assign in2outThrown_payload_endOfPack = videoIn_fork_io_outputs_1_payload_endOfPack;
  always @(*) begin
    feedbackAdded_valid = fifo_pop_fork_io_outputs_0_valid;
    if(feedbackAddCond) begin
      feedbackAdded_valid = 1'b1;
    end
  end

  always @(*) begin
    fifo_pop_fork_io_outputs_0_ready = feedbackAdded_ready;
    if(feedbackAddCond) begin
      fifo_pop_fork_io_outputs_0_ready = 1'b0;
    end
  end

  assign feedbackAdded_payload_0_pixel_0 = fifo_pop_fork_io_outputs_0_payload_0_pixel_0;
  assign feedbackAdded_payload_0_pixel_1 = fifo_pop_fork_io_outputs_0_payload_0_pixel_1;
  assign feedbackAdded_payload_0_pixel_2 = fifo_pop_fork_io_outputs_0_payload_0_pixel_2;
  assign feedbackAdded_payload_0_pixel_3 = fifo_pop_fork_io_outputs_0_payload_0_pixel_3;
  assign feedbackAdded_payload_0_pixel_4 = fifo_pop_fork_io_outputs_0_payload_0_pixel_4;
  assign feedbackAdded_payload_0_pixel_5 = fifo_pop_fork_io_outputs_0_payload_0_pixel_5;
  assign feedbackAdded_payload_0_pixel_6 = fifo_pop_fork_io_outputs_0_payload_0_pixel_6;
  assign feedbackAdded_payload_0_pixel_7 = fifo_pop_fork_io_outputs_0_payload_0_pixel_7;
  assign feedbackAdded_payload_0_pixel_8 = fifo_pop_fork_io_outputs_0_payload_0_pixel_8;
  assign feedbackAdded_payload_0_pixel_9 = fifo_pop_fork_io_outputs_0_payload_0_pixel_9;
  assign feedbackAdded_payload_0_pixel_10 = fifo_pop_fork_io_outputs_0_payload_0_pixel_10;
  assign feedbackAdded_payload_0_pixel_11 = fifo_pop_fork_io_outputs_0_payload_0_pixel_11;
  assign feedbackAdded_payload_0_pixel_12 = fifo_pop_fork_io_outputs_0_payload_0_pixel_12;
  assign feedbackAdded_payload_0_pixel_13 = fifo_pop_fork_io_outputs_0_payload_0_pixel_13;
  assign feedbackAdded_payload_0_pixel_14 = fifo_pop_fork_io_outputs_0_payload_0_pixel_14;
  assign feedbackAdded_payload_0_pixel_15 = fifo_pop_fork_io_outputs_0_payload_0_pixel_15;
  assign feedbackAdded_payload_0_endOfLine = fifo_pop_fork_io_outputs_0_payload_0_endOfLine;
  assign in2fifoJoinFeedback_valid = (videoIn_fork_io_outputs_0_valid && feedbackAdded_valid);
  assign in2fifoJoinFeedback_fire = (in2fifoJoinFeedback_valid && in2fifoJoinFeedback_ready);
  assign in2fifoJoinFeedback_fire_1 = (in2fifoJoinFeedback_valid && in2fifoJoinFeedback_ready);
  assign feedbackAdded_ready = in2fifoJoinFeedback_fire_1;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_0 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_0;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_1 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_1;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_2 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_2;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_3 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_3;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_4 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_4;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_5 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_5;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_6 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_6;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_7 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_7;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_8 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_8;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_9 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_9;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_10 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_10;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_11 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_11;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_12 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_12;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_13 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_13;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_14 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_14;
  assign in2fifoJoinFeedback_payload__1_frame_line_pixel_15 = videoIn_fork_io_outputs_0_payload_frame_line_pixel_15;
  assign in2fifoJoinFeedback_payload__1_frame_line_endOfLine = videoIn_fork_io_outputs_0_payload_frame_line_endOfLine;
  assign in2fifoJoinFeedback_payload__1_frame_endOfFrame = videoIn_fork_io_outputs_0_payload_frame_endOfFrame;
  assign in2fifoJoinFeedback_payload__1_endOfPack = videoIn_fork_io_outputs_0_payload_endOfPack;
  assign in2fifoJoinFeedback_payload__2_0_pixel_0 = feedbackAdded_payload_0_pixel_0;
  assign in2fifoJoinFeedback_payload__2_0_pixel_1 = feedbackAdded_payload_0_pixel_1;
  assign in2fifoJoinFeedback_payload__2_0_pixel_2 = feedbackAdded_payload_0_pixel_2;
  assign in2fifoJoinFeedback_payload__2_0_pixel_3 = feedbackAdded_payload_0_pixel_3;
  assign in2fifoJoinFeedback_payload__2_0_pixel_4 = feedbackAdded_payload_0_pixel_4;
  assign in2fifoJoinFeedback_payload__2_0_pixel_5 = feedbackAdded_payload_0_pixel_5;
  assign in2fifoJoinFeedback_payload__2_0_pixel_6 = feedbackAdded_payload_0_pixel_6;
  assign in2fifoJoinFeedback_payload__2_0_pixel_7 = feedbackAdded_payload_0_pixel_7;
  assign in2fifoJoinFeedback_payload__2_0_pixel_8 = feedbackAdded_payload_0_pixel_8;
  assign in2fifoJoinFeedback_payload__2_0_pixel_9 = feedbackAdded_payload_0_pixel_9;
  assign in2fifoJoinFeedback_payload__2_0_pixel_10 = feedbackAdded_payload_0_pixel_10;
  assign in2fifoJoinFeedback_payload__2_0_pixel_11 = feedbackAdded_payload_0_pixel_11;
  assign in2fifoJoinFeedback_payload__2_0_pixel_12 = feedbackAdded_payload_0_pixel_12;
  assign in2fifoJoinFeedback_payload__2_0_pixel_13 = feedbackAdded_payload_0_pixel_13;
  assign in2fifoJoinFeedback_payload__2_0_pixel_14 = feedbackAdded_payload_0_pixel_14;
  assign in2fifoJoinFeedback_payload__2_0_pixel_15 = feedbackAdded_payload_0_pixel_15;
  assign in2fifoJoinFeedback_payload__2_0_endOfLine = feedbackAdded_payload_0_endOfLine;
  assign in2outJoinFifo2out_valid = (in2outThrown_valid && fifo_pop_fork_io_outputs_1_valid);
  assign in2outJoinFifo2out_fire = (in2outJoinFifo2out_valid && in2outJoinFifo2out_ready);
  assign in2outThrown_ready = in2outJoinFifo2out_fire;
  assign in2outJoinFifo2out_fire_1 = (in2outJoinFifo2out_valid && in2outJoinFifo2out_ready);
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_0 = in2outThrown_payload_frame_line_pixel_0;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_1 = in2outThrown_payload_frame_line_pixel_1;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_2 = in2outThrown_payload_frame_line_pixel_2;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_3 = in2outThrown_payload_frame_line_pixel_3;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_4 = in2outThrown_payload_frame_line_pixel_4;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_5 = in2outThrown_payload_frame_line_pixel_5;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_6 = in2outThrown_payload_frame_line_pixel_6;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_7 = in2outThrown_payload_frame_line_pixel_7;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_8 = in2outThrown_payload_frame_line_pixel_8;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_9 = in2outThrown_payload_frame_line_pixel_9;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_10 = in2outThrown_payload_frame_line_pixel_10;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_11 = in2outThrown_payload_frame_line_pixel_11;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_12 = in2outThrown_payload_frame_line_pixel_12;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_13 = in2outThrown_payload_frame_line_pixel_13;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_14 = in2outThrown_payload_frame_line_pixel_14;
  assign in2outJoinFifo2out_payload__1_frame_line_pixel_15 = in2outThrown_payload_frame_line_pixel_15;
  assign in2outJoinFifo2out_payload__1_frame_line_endOfLine = in2outThrown_payload_frame_line_endOfLine;
  assign in2outJoinFifo2out_payload__1_frame_endOfFrame = in2outThrown_payload_frame_endOfFrame;
  assign in2outJoinFifo2out_payload__1_endOfPack = in2outThrown_payload_endOfPack;
  assign in2outJoinFifo2out_payload__2_0_pixel_0 = fifo_pop_fork_io_outputs_1_payload_0_pixel_0;
  assign in2outJoinFifo2out_payload__2_0_pixel_1 = fifo_pop_fork_io_outputs_1_payload_0_pixel_1;
  assign in2outJoinFifo2out_payload__2_0_pixel_2 = fifo_pop_fork_io_outputs_1_payload_0_pixel_2;
  assign in2outJoinFifo2out_payload__2_0_pixel_3 = fifo_pop_fork_io_outputs_1_payload_0_pixel_3;
  assign in2outJoinFifo2out_payload__2_0_pixel_4 = fifo_pop_fork_io_outputs_1_payload_0_pixel_4;
  assign in2outJoinFifo2out_payload__2_0_pixel_5 = fifo_pop_fork_io_outputs_1_payload_0_pixel_5;
  assign in2outJoinFifo2out_payload__2_0_pixel_6 = fifo_pop_fork_io_outputs_1_payload_0_pixel_6;
  assign in2outJoinFifo2out_payload__2_0_pixel_7 = fifo_pop_fork_io_outputs_1_payload_0_pixel_7;
  assign in2outJoinFifo2out_payload__2_0_pixel_8 = fifo_pop_fork_io_outputs_1_payload_0_pixel_8;
  assign in2outJoinFifo2out_payload__2_0_pixel_9 = fifo_pop_fork_io_outputs_1_payload_0_pixel_9;
  assign in2outJoinFifo2out_payload__2_0_pixel_10 = fifo_pop_fork_io_outputs_1_payload_0_pixel_10;
  assign in2outJoinFifo2out_payload__2_0_pixel_11 = fifo_pop_fork_io_outputs_1_payload_0_pixel_11;
  assign in2outJoinFifo2out_payload__2_0_pixel_12 = fifo_pop_fork_io_outputs_1_payload_0_pixel_12;
  assign in2outJoinFifo2out_payload__2_0_pixel_13 = fifo_pop_fork_io_outputs_1_payload_0_pixel_13;
  assign in2outJoinFifo2out_payload__2_0_pixel_14 = fifo_pop_fork_io_outputs_1_payload_0_pixel_14;
  assign in2outJoinFifo2out_payload__2_0_pixel_15 = fifo_pop_fork_io_outputs_1_payload_0_pixel_15;
  assign in2outJoinFifo2out_payload__2_0_endOfLine = fifo_pop_fork_io_outputs_1_payload_0_endOfLine;
  assign ioVideoInFire = (videoIn_valid && videoIn_ready);
  always @(*) begin
    lineCnt_willIncrement = 1'b0;
    if(when_LineBufferValid_l59) begin
      lineCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    lineCnt_willClear = 1'b0;
    if(when_LineBufferValid_l58) begin
      lineCnt_willClear = 1'b1;
    end
  end

  assign lineCnt_willOverflowIfInc = (lineCnt_value == 1'b1);
  assign lineCnt_willOverflow = (lineCnt_willOverflowIfInc && lineCnt_willIncrement);
  always @(*) begin
    lineCnt_valueNext = (lineCnt_value + lineCnt_willIncrement);
    if(lineCnt_willClear) begin
      lineCnt_valueNext = 1'b0;
    end
  end

  assign lineCntWontOverflowIfInc = (! lineCnt_willOverflowIfInc);
  assign when_LineBufferValid_l58 = (ioVideoInFire && videoIn_payload_frame_endOfFrame);
  assign when_LineBufferValid_l59 = ((ioVideoInFire && videoIn_payload_frame_line_endOfLine) && lineCntWontOverflowIfInc);
  assign in2outThrowCond = lineCntWontOverflowIfInc;
  assign feedbackAddCond = (lineCnt_value == 1'b0);
  assign in2fifoJoinFeedback_ready = fifo_push_ready;
  assign fifo_flush = (ioVideoInFire && videoIn_payload_frame_endOfFrame);
  assign videoOut_valid = in2outJoinFifo2out_valid;
  assign in2outJoinFifo2out_ready = videoOut_ready;
  assign videoOut_payload_endOfPack = videoIn_payload_endOfPack;
  assign videoOut_payload_frame_endOfFrame = videoIn_payload_frame_endOfFrame;
  assign videoOut_payload_frame_line_pixel_0_0 = in2outJoinFifo2out_payload__2_0_pixel_0;
  assign videoOut_payload_frame_line_pixel_0_1 = in2outJoinFifo2out_payload__2_0_pixel_1;
  assign videoOut_payload_frame_line_pixel_0_2 = in2outJoinFifo2out_payload__2_0_pixel_2;
  assign videoOut_payload_frame_line_pixel_0_3 = in2outJoinFifo2out_payload__2_0_pixel_3;
  assign videoOut_payload_frame_line_pixel_0_4 = in2outJoinFifo2out_payload__2_0_pixel_4;
  assign videoOut_payload_frame_line_pixel_0_5 = in2outJoinFifo2out_payload__2_0_pixel_5;
  assign videoOut_payload_frame_line_pixel_0_6 = in2outJoinFifo2out_payload__2_0_pixel_6;
  assign videoOut_payload_frame_line_pixel_0_7 = in2outJoinFifo2out_payload__2_0_pixel_7;
  assign videoOut_payload_frame_line_pixel_0_8 = in2outJoinFifo2out_payload__2_0_pixel_8;
  assign videoOut_payload_frame_line_pixel_0_9 = in2outJoinFifo2out_payload__2_0_pixel_9;
  assign videoOut_payload_frame_line_pixel_0_10 = in2outJoinFifo2out_payload__2_0_pixel_10;
  assign videoOut_payload_frame_line_pixel_0_11 = in2outJoinFifo2out_payload__2_0_pixel_11;
  assign videoOut_payload_frame_line_pixel_0_12 = in2outJoinFifo2out_payload__2_0_pixel_12;
  assign videoOut_payload_frame_line_pixel_0_13 = in2outJoinFifo2out_payload__2_0_pixel_13;
  assign videoOut_payload_frame_line_pixel_0_14 = in2outJoinFifo2out_payload__2_0_pixel_14;
  assign videoOut_payload_frame_line_pixel_0_15 = in2outJoinFifo2out_payload__2_0_pixel_15;
  assign videoOut_payload_frame_line_pixel_1_0 = in2outJoinFifo2out_payload__1_frame_line_pixel_0;
  assign videoOut_payload_frame_line_pixel_1_1 = in2outJoinFifo2out_payload__1_frame_line_pixel_1;
  assign videoOut_payload_frame_line_pixel_1_2 = in2outJoinFifo2out_payload__1_frame_line_pixel_2;
  assign videoOut_payload_frame_line_pixel_1_3 = in2outJoinFifo2out_payload__1_frame_line_pixel_3;
  assign videoOut_payload_frame_line_pixel_1_4 = in2outJoinFifo2out_payload__1_frame_line_pixel_4;
  assign videoOut_payload_frame_line_pixel_1_5 = in2outJoinFifo2out_payload__1_frame_line_pixel_5;
  assign videoOut_payload_frame_line_pixel_1_6 = in2outJoinFifo2out_payload__1_frame_line_pixel_6;
  assign videoOut_payload_frame_line_pixel_1_7 = in2outJoinFifo2out_payload__1_frame_line_pixel_7;
  assign videoOut_payload_frame_line_pixel_1_8 = in2outJoinFifo2out_payload__1_frame_line_pixel_8;
  assign videoOut_payload_frame_line_pixel_1_9 = in2outJoinFifo2out_payload__1_frame_line_pixel_9;
  assign videoOut_payload_frame_line_pixel_1_10 = in2outJoinFifo2out_payload__1_frame_line_pixel_10;
  assign videoOut_payload_frame_line_pixel_1_11 = in2outJoinFifo2out_payload__1_frame_line_pixel_11;
  assign videoOut_payload_frame_line_pixel_1_12 = in2outJoinFifo2out_payload__1_frame_line_pixel_12;
  assign videoOut_payload_frame_line_pixel_1_13 = in2outJoinFifo2out_payload__1_frame_line_pixel_13;
  assign videoOut_payload_frame_line_pixel_1_14 = in2outJoinFifo2out_payload__1_frame_line_pixel_14;
  assign videoOut_payload_frame_line_pixel_1_15 = in2outJoinFifo2out_payload__1_frame_line_pixel_15;
  assign videoOut_payload_frame_line_endOfLine = videoIn_payload_frame_line_endOfLine;
  always @(posedge clk) begin
    if(reset) begin
      lineCnt_value <= 1'b0;
    end else begin
      lineCnt_value <= lineCnt_valueNext;
    end
  end


endmodule

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

//APlusDMultB replaced by APlusDMultB

module APlusDMultB (
  input      [29:0]   A,
  input      [17:0]   B,
  input      [26:0]   D,
  output     [47:0]   P,
  input               CEs_0,
  input               CEs_1,
  input               CEs_2,
  input               CEs_3,
  input               clk
);

  wire       [29:0]   dSP48E2_1_ACOUT;
  wire       [17:0]   dSP48E2_1_BCOUT;
  wire       [47:0]   dSP48E2_1_PCOUT;
  wire       [0:0]    dSP48E2_1_CARRYCASCOUT;
  wire       [0:0]    dSP48E2_1_MULTSIGNOUT;
  wire       [47:0]   dSP48E2_1_P;
  wire       [3:0]    dSP48E2_1_CARRYOUT;
  wire       [7:0]    dSP48E2_1_XOROUT;

  DSP48E2 #(
    .A_INPUT("DIRECT"),
    .B_INPUT("DIRECT"),
    .AMULTSEL("AD"),
    .BMULTSEL("B"),
    .PREADDINSEL("A"),
    .USE_MULT("MULTIPLY"),
    .USE_SIMD("ONE48"),
    .AREG(1),
    .BREG(2),
    .CREG(1),
    .DREG(1),
    .ADREG(1),
    .MREG(1),
    .PREG(1),
    .ACASCREG(1),
    .BCASCREG(1),
    .CARRYINREG(1),
    .CARRYINSELREG(1),
    .INMODEREG(1),
    .OPMODEREG(1),
    .ALUMODEREG(1) 
  ) dSP48E2_1 (
    .CLK              (clk                      ), //i
    .ALUMODE          (4'b0000                  ), //i
    .INMODE           (5'h05                    ), //i
    .OPMODE           (9'h005                   ), //i
    .CARRYINSEL       (3'b000                   ), //i
    .ACIN             (30'h0                    ), //i
    .BCIN             (18'h0                    ), //i
    .PCIN             (48'h0                    ), //i
    .CARRYCASCIN      (1'b0                     ), //i
    .MULTSIGNIN       (1'b0                     ), //i
    .ACOUT            (dSP48E2_1_ACOUT[29:0]    ), //o
    .BCOUT            (dSP48E2_1_BCOUT[17:0]    ), //o
    .PCOUT            (dSP48E2_1_PCOUT[47:0]    ), //o
    .CARRYCASCOUT     (dSP48E2_1_CARRYCASCOUT   ), //o
    .MULTSIGNOUT      (dSP48E2_1_MULTSIGNOUT    ), //o
    .CEA1             (CEs_0                    ), //i
    .CEA2             (1'b0                     ), //i
    .CEB1             (CEs_0                    ), //i
    .CEB2             (CEs_1                    ), //i
    .CEC              (1'b0                     ), //i
    .CED              (CEs_0                    ), //i
    .CEAD             (CEs_1                    ), //i
    .CEM              (CEs_2                    ), //i
    .CEP              (CEs_3                    ), //i
    .CECARRYIN        (1'b0                     ), //i
    .CECTRL           (1'b0                     ), //i
    .CEINMODE         (1'b0                     ), //i
    .CEALUMODE        (1'b0                     ), //i
    .RSTA             (1'b0                     ), //i
    .RSTB             (1'b0                     ), //i
    .RSTC             (1'b0                     ), //i
    .RSTD             (1'b0                     ), //i
    .RSTM             (1'b0                     ), //i
    .RSTP             (1'b0                     ), //i
    .RSTALLCARRYIN    (1'b0                     ), //i
    .RSTCTRL          (1'b0                     ), //i
    .RSTINMODE        (1'b0                     ), //i
    .RSTALUMODE       (1'b0                     ), //i
    .A                (A[29:0]                  ), //i
    .B                (B[17:0]                  ), //i
    .C                (48'h0                    ), //i
    .D                (D[26:0]                  ), //i
    .CARRYIN          (1'b0                     ), //i
    .P                (dSP48E2_1_P[47:0]        ), //o
    .CARRYOUT         (dSP48E2_1_CARRYOUT[3:0]  ), //o
    .XOROUT           (dSP48E2_1_XOROUT[7:0]    )  //o
  );
  assign P = dSP48E2_1_P;

endmodule

module StreamFork_3 (
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_0_pixel_0,
  input      [7:0]    io_input_payload_0_pixel_1,
  input      [7:0]    io_input_payload_0_pixel_2,
  input      [7:0]    io_input_payload_0_pixel_3,
  input      [7:0]    io_input_payload_0_pixel_4,
  input      [7:0]    io_input_payload_0_pixel_5,
  input      [7:0]    io_input_payload_0_pixel_6,
  input      [7:0]    io_input_payload_0_pixel_7,
  input      [7:0]    io_input_payload_0_pixel_8,
  input      [7:0]    io_input_payload_0_pixel_9,
  input      [7:0]    io_input_payload_0_pixel_10,
  input      [7:0]    io_input_payload_0_pixel_11,
  input      [7:0]    io_input_payload_0_pixel_12,
  input      [7:0]    io_input_payload_0_pixel_13,
  input      [7:0]    io_input_payload_0_pixel_14,
  input      [7:0]    io_input_payload_0_pixel_15,
  input               io_input_payload_0_endOfLine,
  input      [7:0]    io_input_payload_1_pixel_0,
  input      [7:0]    io_input_payload_1_pixel_1,
  input      [7:0]    io_input_payload_1_pixel_2,
  input      [7:0]    io_input_payload_1_pixel_3,
  input      [7:0]    io_input_payload_1_pixel_4,
  input      [7:0]    io_input_payload_1_pixel_5,
  input      [7:0]    io_input_payload_1_pixel_6,
  input      [7:0]    io_input_payload_1_pixel_7,
  input      [7:0]    io_input_payload_1_pixel_8,
  input      [7:0]    io_input_payload_1_pixel_9,
  input      [7:0]    io_input_payload_1_pixel_10,
  input      [7:0]    io_input_payload_1_pixel_11,
  input      [7:0]    io_input_payload_1_pixel_12,
  input      [7:0]    io_input_payload_1_pixel_13,
  input      [7:0]    io_input_payload_1_pixel_14,
  input      [7:0]    io_input_payload_1_pixel_15,
  input               io_input_payload_1_endOfLine,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_0_pixel_0,
  output     [7:0]    io_outputs_0_payload_0_pixel_1,
  output     [7:0]    io_outputs_0_payload_0_pixel_2,
  output     [7:0]    io_outputs_0_payload_0_pixel_3,
  output     [7:0]    io_outputs_0_payload_0_pixel_4,
  output     [7:0]    io_outputs_0_payload_0_pixel_5,
  output     [7:0]    io_outputs_0_payload_0_pixel_6,
  output     [7:0]    io_outputs_0_payload_0_pixel_7,
  output     [7:0]    io_outputs_0_payload_0_pixel_8,
  output     [7:0]    io_outputs_0_payload_0_pixel_9,
  output     [7:0]    io_outputs_0_payload_0_pixel_10,
  output     [7:0]    io_outputs_0_payload_0_pixel_11,
  output     [7:0]    io_outputs_0_payload_0_pixel_12,
  output     [7:0]    io_outputs_0_payload_0_pixel_13,
  output     [7:0]    io_outputs_0_payload_0_pixel_14,
  output     [7:0]    io_outputs_0_payload_0_pixel_15,
  output              io_outputs_0_payload_0_endOfLine,
  output     [7:0]    io_outputs_0_payload_1_pixel_0,
  output     [7:0]    io_outputs_0_payload_1_pixel_1,
  output     [7:0]    io_outputs_0_payload_1_pixel_2,
  output     [7:0]    io_outputs_0_payload_1_pixel_3,
  output     [7:0]    io_outputs_0_payload_1_pixel_4,
  output     [7:0]    io_outputs_0_payload_1_pixel_5,
  output     [7:0]    io_outputs_0_payload_1_pixel_6,
  output     [7:0]    io_outputs_0_payload_1_pixel_7,
  output     [7:0]    io_outputs_0_payload_1_pixel_8,
  output     [7:0]    io_outputs_0_payload_1_pixel_9,
  output     [7:0]    io_outputs_0_payload_1_pixel_10,
  output     [7:0]    io_outputs_0_payload_1_pixel_11,
  output     [7:0]    io_outputs_0_payload_1_pixel_12,
  output     [7:0]    io_outputs_0_payload_1_pixel_13,
  output     [7:0]    io_outputs_0_payload_1_pixel_14,
  output     [7:0]    io_outputs_0_payload_1_pixel_15,
  output              io_outputs_0_payload_1_endOfLine,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_0_pixel_0,
  output     [7:0]    io_outputs_1_payload_0_pixel_1,
  output     [7:0]    io_outputs_1_payload_0_pixel_2,
  output     [7:0]    io_outputs_1_payload_0_pixel_3,
  output     [7:0]    io_outputs_1_payload_0_pixel_4,
  output     [7:0]    io_outputs_1_payload_0_pixel_5,
  output     [7:0]    io_outputs_1_payload_0_pixel_6,
  output     [7:0]    io_outputs_1_payload_0_pixel_7,
  output     [7:0]    io_outputs_1_payload_0_pixel_8,
  output     [7:0]    io_outputs_1_payload_0_pixel_9,
  output     [7:0]    io_outputs_1_payload_0_pixel_10,
  output     [7:0]    io_outputs_1_payload_0_pixel_11,
  output     [7:0]    io_outputs_1_payload_0_pixel_12,
  output     [7:0]    io_outputs_1_payload_0_pixel_13,
  output     [7:0]    io_outputs_1_payload_0_pixel_14,
  output     [7:0]    io_outputs_1_payload_0_pixel_15,
  output              io_outputs_1_payload_0_endOfLine,
  output     [7:0]    io_outputs_1_payload_1_pixel_0,
  output     [7:0]    io_outputs_1_payload_1_pixel_1,
  output     [7:0]    io_outputs_1_payload_1_pixel_2,
  output     [7:0]    io_outputs_1_payload_1_pixel_3,
  output     [7:0]    io_outputs_1_payload_1_pixel_4,
  output     [7:0]    io_outputs_1_payload_1_pixel_5,
  output     [7:0]    io_outputs_1_payload_1_pixel_6,
  output     [7:0]    io_outputs_1_payload_1_pixel_7,
  output     [7:0]    io_outputs_1_payload_1_pixel_8,
  output     [7:0]    io_outputs_1_payload_1_pixel_9,
  output     [7:0]    io_outputs_1_payload_1_pixel_10,
  output     [7:0]    io_outputs_1_payload_1_pixel_11,
  output     [7:0]    io_outputs_1_payload_1_pixel_12,
  output     [7:0]    io_outputs_1_payload_1_pixel_13,
  output     [7:0]    io_outputs_1_payload_1_pixel_14,
  output     [7:0]    io_outputs_1_payload_1_pixel_15,
  output              io_outputs_1_payload_1_endOfLine,
  input               clk,
  input               reset
);

  reg                 tmp_io_outputs_0_valid;
  reg                 tmp_io_outputs_1_valid;
  wire                when_Stream_l825;
  wire                when_Stream_l825_1;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l825) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_1) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l825 = ((! io_outputs_0_ready) && tmp_io_outputs_0_valid);
  assign when_Stream_l825_1 = ((! io_outputs_1_ready) && tmp_io_outputs_1_valid);
  assign io_outputs_0_valid = (io_input_valid && tmp_io_outputs_0_valid);
  assign io_outputs_0_payload_0_pixel_0 = io_input_payload_0_pixel_0;
  assign io_outputs_0_payload_0_pixel_1 = io_input_payload_0_pixel_1;
  assign io_outputs_0_payload_0_pixel_2 = io_input_payload_0_pixel_2;
  assign io_outputs_0_payload_0_pixel_3 = io_input_payload_0_pixel_3;
  assign io_outputs_0_payload_0_pixel_4 = io_input_payload_0_pixel_4;
  assign io_outputs_0_payload_0_pixel_5 = io_input_payload_0_pixel_5;
  assign io_outputs_0_payload_0_pixel_6 = io_input_payload_0_pixel_6;
  assign io_outputs_0_payload_0_pixel_7 = io_input_payload_0_pixel_7;
  assign io_outputs_0_payload_0_pixel_8 = io_input_payload_0_pixel_8;
  assign io_outputs_0_payload_0_pixel_9 = io_input_payload_0_pixel_9;
  assign io_outputs_0_payload_0_pixel_10 = io_input_payload_0_pixel_10;
  assign io_outputs_0_payload_0_pixel_11 = io_input_payload_0_pixel_11;
  assign io_outputs_0_payload_0_pixel_12 = io_input_payload_0_pixel_12;
  assign io_outputs_0_payload_0_pixel_13 = io_input_payload_0_pixel_13;
  assign io_outputs_0_payload_0_pixel_14 = io_input_payload_0_pixel_14;
  assign io_outputs_0_payload_0_pixel_15 = io_input_payload_0_pixel_15;
  assign io_outputs_0_payload_0_endOfLine = io_input_payload_0_endOfLine;
  assign io_outputs_0_payload_1_pixel_0 = io_input_payload_1_pixel_0;
  assign io_outputs_0_payload_1_pixel_1 = io_input_payload_1_pixel_1;
  assign io_outputs_0_payload_1_pixel_2 = io_input_payload_1_pixel_2;
  assign io_outputs_0_payload_1_pixel_3 = io_input_payload_1_pixel_3;
  assign io_outputs_0_payload_1_pixel_4 = io_input_payload_1_pixel_4;
  assign io_outputs_0_payload_1_pixel_5 = io_input_payload_1_pixel_5;
  assign io_outputs_0_payload_1_pixel_6 = io_input_payload_1_pixel_6;
  assign io_outputs_0_payload_1_pixel_7 = io_input_payload_1_pixel_7;
  assign io_outputs_0_payload_1_pixel_8 = io_input_payload_1_pixel_8;
  assign io_outputs_0_payload_1_pixel_9 = io_input_payload_1_pixel_9;
  assign io_outputs_0_payload_1_pixel_10 = io_input_payload_1_pixel_10;
  assign io_outputs_0_payload_1_pixel_11 = io_input_payload_1_pixel_11;
  assign io_outputs_0_payload_1_pixel_12 = io_input_payload_1_pixel_12;
  assign io_outputs_0_payload_1_pixel_13 = io_input_payload_1_pixel_13;
  assign io_outputs_0_payload_1_pixel_14 = io_input_payload_1_pixel_14;
  assign io_outputs_0_payload_1_pixel_15 = io_input_payload_1_pixel_15;
  assign io_outputs_0_payload_1_endOfLine = io_input_payload_1_endOfLine;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && tmp_io_outputs_1_valid);
  assign io_outputs_1_payload_0_pixel_0 = io_input_payload_0_pixel_0;
  assign io_outputs_1_payload_0_pixel_1 = io_input_payload_0_pixel_1;
  assign io_outputs_1_payload_0_pixel_2 = io_input_payload_0_pixel_2;
  assign io_outputs_1_payload_0_pixel_3 = io_input_payload_0_pixel_3;
  assign io_outputs_1_payload_0_pixel_4 = io_input_payload_0_pixel_4;
  assign io_outputs_1_payload_0_pixel_5 = io_input_payload_0_pixel_5;
  assign io_outputs_1_payload_0_pixel_6 = io_input_payload_0_pixel_6;
  assign io_outputs_1_payload_0_pixel_7 = io_input_payload_0_pixel_7;
  assign io_outputs_1_payload_0_pixel_8 = io_input_payload_0_pixel_8;
  assign io_outputs_1_payload_0_pixel_9 = io_input_payload_0_pixel_9;
  assign io_outputs_1_payload_0_pixel_10 = io_input_payload_0_pixel_10;
  assign io_outputs_1_payload_0_pixel_11 = io_input_payload_0_pixel_11;
  assign io_outputs_1_payload_0_pixel_12 = io_input_payload_0_pixel_12;
  assign io_outputs_1_payload_0_pixel_13 = io_input_payload_0_pixel_13;
  assign io_outputs_1_payload_0_pixel_14 = io_input_payload_0_pixel_14;
  assign io_outputs_1_payload_0_pixel_15 = io_input_payload_0_pixel_15;
  assign io_outputs_1_payload_0_endOfLine = io_input_payload_0_endOfLine;
  assign io_outputs_1_payload_1_pixel_0 = io_input_payload_1_pixel_0;
  assign io_outputs_1_payload_1_pixel_1 = io_input_payload_1_pixel_1;
  assign io_outputs_1_payload_1_pixel_2 = io_input_payload_1_pixel_2;
  assign io_outputs_1_payload_1_pixel_3 = io_input_payload_1_pixel_3;
  assign io_outputs_1_payload_1_pixel_4 = io_input_payload_1_pixel_4;
  assign io_outputs_1_payload_1_pixel_5 = io_input_payload_1_pixel_5;
  assign io_outputs_1_payload_1_pixel_6 = io_input_payload_1_pixel_6;
  assign io_outputs_1_payload_1_pixel_7 = io_input_payload_1_pixel_7;
  assign io_outputs_1_payload_1_pixel_8 = io_input_payload_1_pixel_8;
  assign io_outputs_1_payload_1_pixel_9 = io_input_payload_1_pixel_9;
  assign io_outputs_1_payload_1_pixel_10 = io_input_payload_1_pixel_10;
  assign io_outputs_1_payload_1_pixel_11 = io_input_payload_1_pixel_11;
  assign io_outputs_1_payload_1_pixel_12 = io_input_payload_1_pixel_12;
  assign io_outputs_1_payload_1_pixel_13 = io_input_payload_1_pixel_13;
  assign io_outputs_1_payload_1_pixel_14 = io_input_payload_1_pixel_14;
  assign io_outputs_1_payload_1_pixel_15 = io_input_payload_1_pixel_15;
  assign io_outputs_1_payload_1_endOfLine = io_input_payload_1_endOfLine;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  always @(posedge clk) begin
    if(reset) begin
      tmp_io_outputs_0_valid <= 1'b1;
      tmp_io_outputs_1_valid <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        tmp_io_outputs_0_valid <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        tmp_io_outputs_1_valid <= 1'b0;
      end
      if(io_input_ready) begin
        tmp_io_outputs_0_valid <= 1'b1;
        tmp_io_outputs_1_valid <= 1'b1;
      end
    end
  end


endmodule

//StreamFork replaced by StreamFork

module StreamFifoHighPerf_1 (
  input               push_valid,
  output              push_ready,
  input      [7:0]    push_payload_0_pixel_0,
  input      [7:0]    push_payload_0_pixel_1,
  input      [7:0]    push_payload_0_pixel_2,
  input      [7:0]    push_payload_0_pixel_3,
  input      [7:0]    push_payload_0_pixel_4,
  input      [7:0]    push_payload_0_pixel_5,
  input      [7:0]    push_payload_0_pixel_6,
  input      [7:0]    push_payload_0_pixel_7,
  input      [7:0]    push_payload_0_pixel_8,
  input      [7:0]    push_payload_0_pixel_9,
  input      [7:0]    push_payload_0_pixel_10,
  input      [7:0]    push_payload_0_pixel_11,
  input      [7:0]    push_payload_0_pixel_12,
  input      [7:0]    push_payload_0_pixel_13,
  input      [7:0]    push_payload_0_pixel_14,
  input      [7:0]    push_payload_0_pixel_15,
  input               push_payload_0_endOfLine,
  input      [7:0]    push_payload_1_pixel_0,
  input      [7:0]    push_payload_1_pixel_1,
  input      [7:0]    push_payload_1_pixel_2,
  input      [7:0]    push_payload_1_pixel_3,
  input      [7:0]    push_payload_1_pixel_4,
  input      [7:0]    push_payload_1_pixel_5,
  input      [7:0]    push_payload_1_pixel_6,
  input      [7:0]    push_payload_1_pixel_7,
  input      [7:0]    push_payload_1_pixel_8,
  input      [7:0]    push_payload_1_pixel_9,
  input      [7:0]    push_payload_1_pixel_10,
  input      [7:0]    push_payload_1_pixel_11,
  input      [7:0]    push_payload_1_pixel_12,
  input      [7:0]    push_payload_1_pixel_13,
  input      [7:0]    push_payload_1_pixel_14,
  input      [7:0]    push_payload_1_pixel_15,
  input               push_payload_1_endOfLine,
  output              pop_valid,
  input               pop_ready,
  output     [7:0]    pop_payload_0_pixel_0,
  output     [7:0]    pop_payload_0_pixel_1,
  output     [7:0]    pop_payload_0_pixel_2,
  output     [7:0]    pop_payload_0_pixel_3,
  output     [7:0]    pop_payload_0_pixel_4,
  output     [7:0]    pop_payload_0_pixel_5,
  output     [7:0]    pop_payload_0_pixel_6,
  output     [7:0]    pop_payload_0_pixel_7,
  output     [7:0]    pop_payload_0_pixel_8,
  output     [7:0]    pop_payload_0_pixel_9,
  output     [7:0]    pop_payload_0_pixel_10,
  output     [7:0]    pop_payload_0_pixel_11,
  output     [7:0]    pop_payload_0_pixel_12,
  output     [7:0]    pop_payload_0_pixel_13,
  output     [7:0]    pop_payload_0_pixel_14,
  output     [7:0]    pop_payload_0_pixel_15,
  output              pop_payload_0_endOfLine,
  output     [7:0]    pop_payload_1_pixel_0,
  output     [7:0]    pop_payload_1_pixel_1,
  output     [7:0]    pop_payload_1_pixel_2,
  output     [7:0]    pop_payload_1_pixel_3,
  output     [7:0]    pop_payload_1_pixel_4,
  output     [7:0]    pop_payload_1_pixel_5,
  output     [7:0]    pop_payload_1_pixel_6,
  output     [7:0]    pop_payload_1_pixel_7,
  output     [7:0]    pop_payload_1_pixel_8,
  output     [7:0]    pop_payload_1_pixel_9,
  output     [7:0]    pop_payload_1_pixel_10,
  output     [7:0]    pop_payload_1_pixel_11,
  output     [7:0]    pop_payload_1_pixel_12,
  output     [7:0]    pop_payload_1_pixel_13,
  output     [7:0]    pop_payload_1_pixel_14,
  output     [7:0]    pop_payload_1_pixel_15,
  output              pop_payload_1_endOfLine,
  input               flush,
  input               clk,
  input               reset
);

  reg        [257:0]  tmp_ram_port0;
  wire       [8:0]    tmp_pushPtr_valueNext;
  wire       [0:0]    tmp_pushPtr_valueNext_1;
  wire       [8:0]    tmp_popPtr_valueNext;
  wire       [0:0]    tmp_popPtr_valueNext_1;
  wire       [257:0]  tmp_ram_port;
  reg                 tmp_1;
  wire                popEvent_valid;
  reg                 popEvent_ready;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [8:0]    pushPtr_valueNext;
  reg        [8:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [8:0]    popPtr_valueNext;
  reg        [8:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                pushing;
  wire                popping;
  wire                empty;
  wire                full;
  reg                 tmp_popEvent_valid;
  reg                 rValid;
  wire       [7:0]    rData_0_pixel_0;
  wire       [7:0]    rData_0_pixel_1;
  wire       [7:0]    rData_0_pixel_2;
  wire       [7:0]    rData_0_pixel_3;
  wire       [7:0]    rData_0_pixel_4;
  wire       [7:0]    rData_0_pixel_5;
  wire       [7:0]    rData_0_pixel_6;
  wire       [7:0]    rData_0_pixel_7;
  wire       [7:0]    rData_0_pixel_8;
  wire       [7:0]    rData_0_pixel_9;
  wire       [7:0]    rData_0_pixel_10;
  wire       [7:0]    rData_0_pixel_11;
  wire       [7:0]    rData_0_pixel_12;
  wire       [7:0]    rData_0_pixel_13;
  wire       [7:0]    rData_0_pixel_14;
  wire       [7:0]    rData_0_pixel_15;
  wire                rData_0_endOfLine;
  wire       [7:0]    rData_1_pixel_0;
  wire       [7:0]    rData_1_pixel_1;
  wire       [7:0]    rData_1_pixel_2;
  wire       [7:0]    rData_1_pixel_3;
  wire       [7:0]    rData_1_pixel_4;
  wire       [7:0]    rData_1_pixel_5;
  wire       [7:0]    rData_1_pixel_6;
  wire       [7:0]    rData_1_pixel_7;
  wire       [7:0]    rData_1_pixel_8;
  wire       [7:0]    rData_1_pixel_9;
  wire       [7:0]    rData_1_pixel_10;
  wire       [7:0]    rData_1_pixel_11;
  wire       [7:0]    rData_1_pixel_12;
  wire       [7:0]    rData_1_pixel_13;
  wire       [7:0]    rData_1_pixel_14;
  wire       [7:0]    rData_1_pixel_15;
  wire                rData_1_endOfLine;
  wire       [257:0]  tmp_rData_0_pixel_0;
  wire       [128:0]  tmp_rData_0_pixel_0_1;
  wire       [127:0]  tmp_rData_0_pixel_0_2;
  wire       [128:0]  tmp_rData_1_pixel_0;
  wire       [127:0]  tmp_rData_1_pixel_0_1;
  wire                when_StreamFifoHighPerf_l38;
  wire                when_StreamFifoHighPerf_l42;
  reg [257:0] ram [0:511];

  assign tmp_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign tmp_pushPtr_valueNext = {8'd0, tmp_pushPtr_valueNext_1};
  assign tmp_popPtr_valueNext_1 = popPtr_willIncrement;
  assign tmp_popPtr_valueNext = {8'd0, tmp_popPtr_valueNext_1};
  assign tmp_ram_port = {{push_payload_1_endOfLine,{push_payload_1_pixel_15,{push_payload_1_pixel_14,{push_payload_1_pixel_13,{push_payload_1_pixel_12,{push_payload_1_pixel_11,{push_payload_1_pixel_10,{push_payload_1_pixel_9,{push_payload_1_pixel_8,{push_payload_1_pixel_7,{push_payload_1_pixel_6,{push_payload_1_pixel_5,{push_payload_1_pixel_4,{push_payload_1_pixel_3,{push_payload_1_pixel_2,{push_payload_1_pixel_1,push_payload_1_pixel_0}}}}}}}}}}}}}}}},{push_payload_0_endOfLine,{push_payload_0_pixel_15,{push_payload_0_pixel_14,{push_payload_0_pixel_13,{push_payload_0_pixel_12,{push_payload_0_pixel_11,{push_payload_0_pixel_10,{push_payload_0_pixel_9,{push_payload_0_pixel_8,{push_payload_0_pixel_7,{push_payload_0_pixel_6,{push_payload_0_pixel_5,{push_payload_0_pixel_4,{push_payload_0_pixel_3,{push_payload_0_pixel_2,{push_payload_0_pixel_1,push_payload_0_pixel_0}}}}}}}}}}}}}}}}};
  always @(posedge clk) begin
    if(popEvent_ready) begin
      tmp_ram_port0 <= ram[popPtr_value];
    end
  end

  always @(posedge clk) begin
    if(tmp_1) begin
      ram[pushPtr_value] <= tmp_ram_port;
    end
  end

  always @(*) begin
    tmp_1 = 1'b0;
    if(pushing) begin
      tmp_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 9'h1ff);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + tmp_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 9'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 9'h1ff);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + tmp_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 9'h0;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign pushing = (push_valid && push_ready);
  assign popping = (popEvent_valid && popEvent_ready);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign push_ready = (! full);
  assign popEvent_valid = ((! empty) && (! (tmp_popEvent_valid && (! full))));
  assign tmp_rData_0_pixel_0 = tmp_ram_port0;
  assign tmp_rData_0_pixel_0_1 = tmp_rData_0_pixel_0[128 : 0];
  assign tmp_rData_0_pixel_0_2 = tmp_rData_0_pixel_0_1[127 : 0];
  assign rData_0_pixel_0 = tmp_rData_0_pixel_0_2[7 : 0];
  assign rData_0_pixel_1 = tmp_rData_0_pixel_0_2[15 : 8];
  assign rData_0_pixel_2 = tmp_rData_0_pixel_0_2[23 : 16];
  assign rData_0_pixel_3 = tmp_rData_0_pixel_0_2[31 : 24];
  assign rData_0_pixel_4 = tmp_rData_0_pixel_0_2[39 : 32];
  assign rData_0_pixel_5 = tmp_rData_0_pixel_0_2[47 : 40];
  assign rData_0_pixel_6 = tmp_rData_0_pixel_0_2[55 : 48];
  assign rData_0_pixel_7 = tmp_rData_0_pixel_0_2[63 : 56];
  assign rData_0_pixel_8 = tmp_rData_0_pixel_0_2[71 : 64];
  assign rData_0_pixel_9 = tmp_rData_0_pixel_0_2[79 : 72];
  assign rData_0_pixel_10 = tmp_rData_0_pixel_0_2[87 : 80];
  assign rData_0_pixel_11 = tmp_rData_0_pixel_0_2[95 : 88];
  assign rData_0_pixel_12 = tmp_rData_0_pixel_0_2[103 : 96];
  assign rData_0_pixel_13 = tmp_rData_0_pixel_0_2[111 : 104];
  assign rData_0_pixel_14 = tmp_rData_0_pixel_0_2[119 : 112];
  assign rData_0_pixel_15 = tmp_rData_0_pixel_0_2[127 : 120];
  assign rData_0_endOfLine = tmp_rData_0_pixel_0_1[128];
  assign tmp_rData_1_pixel_0 = tmp_rData_0_pixel_0[257 : 129];
  assign tmp_rData_1_pixel_0_1 = tmp_rData_1_pixel_0[127 : 0];
  assign rData_1_pixel_0 = tmp_rData_1_pixel_0_1[7 : 0];
  assign rData_1_pixel_1 = tmp_rData_1_pixel_0_1[15 : 8];
  assign rData_1_pixel_2 = tmp_rData_1_pixel_0_1[23 : 16];
  assign rData_1_pixel_3 = tmp_rData_1_pixel_0_1[31 : 24];
  assign rData_1_pixel_4 = tmp_rData_1_pixel_0_1[39 : 32];
  assign rData_1_pixel_5 = tmp_rData_1_pixel_0_1[47 : 40];
  assign rData_1_pixel_6 = tmp_rData_1_pixel_0_1[55 : 48];
  assign rData_1_pixel_7 = tmp_rData_1_pixel_0_1[63 : 56];
  assign rData_1_pixel_8 = tmp_rData_1_pixel_0_1[71 : 64];
  assign rData_1_pixel_9 = tmp_rData_1_pixel_0_1[79 : 72];
  assign rData_1_pixel_10 = tmp_rData_1_pixel_0_1[87 : 80];
  assign rData_1_pixel_11 = tmp_rData_1_pixel_0_1[95 : 88];
  assign rData_1_pixel_12 = tmp_rData_1_pixel_0_1[103 : 96];
  assign rData_1_pixel_13 = tmp_rData_1_pixel_0_1[111 : 104];
  assign rData_1_pixel_14 = tmp_rData_1_pixel_0_1[119 : 112];
  assign rData_1_pixel_15 = tmp_rData_1_pixel_0_1[127 : 120];
  assign rData_1_endOfLine = tmp_rData_1_pixel_0[128];
  always @(*) begin
    popEvent_ready = pop_ready;
    if(when_StreamFifoHighPerf_l38) begin
      popEvent_ready = 1'b1;
    end
  end

  assign when_StreamFifoHighPerf_l38 = (! rValid);
  assign pop_valid = rValid;
  assign pop_payload_0_pixel_0 = rData_0_pixel_0;
  assign pop_payload_0_pixel_1 = rData_0_pixel_1;
  assign pop_payload_0_pixel_2 = rData_0_pixel_2;
  assign pop_payload_0_pixel_3 = rData_0_pixel_3;
  assign pop_payload_0_pixel_4 = rData_0_pixel_4;
  assign pop_payload_0_pixel_5 = rData_0_pixel_5;
  assign pop_payload_0_pixel_6 = rData_0_pixel_6;
  assign pop_payload_0_pixel_7 = rData_0_pixel_7;
  assign pop_payload_0_pixel_8 = rData_0_pixel_8;
  assign pop_payload_0_pixel_9 = rData_0_pixel_9;
  assign pop_payload_0_pixel_10 = rData_0_pixel_10;
  assign pop_payload_0_pixel_11 = rData_0_pixel_11;
  assign pop_payload_0_pixel_12 = rData_0_pixel_12;
  assign pop_payload_0_pixel_13 = rData_0_pixel_13;
  assign pop_payload_0_pixel_14 = rData_0_pixel_14;
  assign pop_payload_0_pixel_15 = rData_0_pixel_15;
  assign pop_payload_0_endOfLine = rData_0_endOfLine;
  assign pop_payload_1_pixel_0 = rData_1_pixel_0;
  assign pop_payload_1_pixel_1 = rData_1_pixel_1;
  assign pop_payload_1_pixel_2 = rData_1_pixel_2;
  assign pop_payload_1_pixel_3 = rData_1_pixel_3;
  assign pop_payload_1_pixel_4 = rData_1_pixel_4;
  assign pop_payload_1_pixel_5 = rData_1_pixel_5;
  assign pop_payload_1_pixel_6 = rData_1_pixel_6;
  assign pop_payload_1_pixel_7 = rData_1_pixel_7;
  assign pop_payload_1_pixel_8 = rData_1_pixel_8;
  assign pop_payload_1_pixel_9 = rData_1_pixel_9;
  assign pop_payload_1_pixel_10 = rData_1_pixel_10;
  assign pop_payload_1_pixel_11 = rData_1_pixel_11;
  assign pop_payload_1_pixel_12 = rData_1_pixel_12;
  assign pop_payload_1_pixel_13 = rData_1_pixel_13;
  assign pop_payload_1_pixel_14 = rData_1_pixel_14;
  assign pop_payload_1_pixel_15 = rData_1_pixel_15;
  assign pop_payload_1_endOfLine = rData_1_endOfLine;
  assign when_StreamFifoHighPerf_l42 = (pushing != popping);
  always @(posedge clk) begin
    if(reset) begin
      pushPtr_value <= 9'h0;
      popPtr_value <= 9'h0;
      risingOccupancy <= 1'b0;
      tmp_popEvent_valid <= 1'b0;
      rValid <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      tmp_popEvent_valid <= (popPtr_valueNext == pushPtr_value);
      if(popEvent_ready) begin
        rValid <= popEvent_valid;
      end
      if(when_StreamFifoHighPerf_l42) begin
        risingOccupancy <= pushing;
      end
      if(flush) begin
        rValid <= 1'b0;
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamFork_1 (
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_0_pixel_0,
  input      [7:0]    io_input_payload_0_pixel_1,
  input      [7:0]    io_input_payload_0_pixel_2,
  input      [7:0]    io_input_payload_0_pixel_3,
  input      [7:0]    io_input_payload_0_pixel_4,
  input      [7:0]    io_input_payload_0_pixel_5,
  input      [7:0]    io_input_payload_0_pixel_6,
  input      [7:0]    io_input_payload_0_pixel_7,
  input      [7:0]    io_input_payload_0_pixel_8,
  input      [7:0]    io_input_payload_0_pixel_9,
  input      [7:0]    io_input_payload_0_pixel_10,
  input      [7:0]    io_input_payload_0_pixel_11,
  input      [7:0]    io_input_payload_0_pixel_12,
  input      [7:0]    io_input_payload_0_pixel_13,
  input      [7:0]    io_input_payload_0_pixel_14,
  input      [7:0]    io_input_payload_0_pixel_15,
  input               io_input_payload_0_endOfLine,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_0_pixel_0,
  output     [7:0]    io_outputs_0_payload_0_pixel_1,
  output     [7:0]    io_outputs_0_payload_0_pixel_2,
  output     [7:0]    io_outputs_0_payload_0_pixel_3,
  output     [7:0]    io_outputs_0_payload_0_pixel_4,
  output     [7:0]    io_outputs_0_payload_0_pixel_5,
  output     [7:0]    io_outputs_0_payload_0_pixel_6,
  output     [7:0]    io_outputs_0_payload_0_pixel_7,
  output     [7:0]    io_outputs_0_payload_0_pixel_8,
  output     [7:0]    io_outputs_0_payload_0_pixel_9,
  output     [7:0]    io_outputs_0_payload_0_pixel_10,
  output     [7:0]    io_outputs_0_payload_0_pixel_11,
  output     [7:0]    io_outputs_0_payload_0_pixel_12,
  output     [7:0]    io_outputs_0_payload_0_pixel_13,
  output     [7:0]    io_outputs_0_payload_0_pixel_14,
  output     [7:0]    io_outputs_0_payload_0_pixel_15,
  output              io_outputs_0_payload_0_endOfLine,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_0_pixel_0,
  output     [7:0]    io_outputs_1_payload_0_pixel_1,
  output     [7:0]    io_outputs_1_payload_0_pixel_2,
  output     [7:0]    io_outputs_1_payload_0_pixel_3,
  output     [7:0]    io_outputs_1_payload_0_pixel_4,
  output     [7:0]    io_outputs_1_payload_0_pixel_5,
  output     [7:0]    io_outputs_1_payload_0_pixel_6,
  output     [7:0]    io_outputs_1_payload_0_pixel_7,
  output     [7:0]    io_outputs_1_payload_0_pixel_8,
  output     [7:0]    io_outputs_1_payload_0_pixel_9,
  output     [7:0]    io_outputs_1_payload_0_pixel_10,
  output     [7:0]    io_outputs_1_payload_0_pixel_11,
  output     [7:0]    io_outputs_1_payload_0_pixel_12,
  output     [7:0]    io_outputs_1_payload_0_pixel_13,
  output     [7:0]    io_outputs_1_payload_0_pixel_14,
  output     [7:0]    io_outputs_1_payload_0_pixel_15,
  output              io_outputs_1_payload_0_endOfLine,
  input               clk,
  input               reset
);

  reg                 tmp_io_outputs_0_valid;
  reg                 tmp_io_outputs_1_valid;
  wire                when_Stream_l825;
  wire                when_Stream_l825_1;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l825) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_1) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l825 = ((! io_outputs_0_ready) && tmp_io_outputs_0_valid);
  assign when_Stream_l825_1 = ((! io_outputs_1_ready) && tmp_io_outputs_1_valid);
  assign io_outputs_0_valid = (io_input_valid && tmp_io_outputs_0_valid);
  assign io_outputs_0_payload_0_pixel_0 = io_input_payload_0_pixel_0;
  assign io_outputs_0_payload_0_pixel_1 = io_input_payload_0_pixel_1;
  assign io_outputs_0_payload_0_pixel_2 = io_input_payload_0_pixel_2;
  assign io_outputs_0_payload_0_pixel_3 = io_input_payload_0_pixel_3;
  assign io_outputs_0_payload_0_pixel_4 = io_input_payload_0_pixel_4;
  assign io_outputs_0_payload_0_pixel_5 = io_input_payload_0_pixel_5;
  assign io_outputs_0_payload_0_pixel_6 = io_input_payload_0_pixel_6;
  assign io_outputs_0_payload_0_pixel_7 = io_input_payload_0_pixel_7;
  assign io_outputs_0_payload_0_pixel_8 = io_input_payload_0_pixel_8;
  assign io_outputs_0_payload_0_pixel_9 = io_input_payload_0_pixel_9;
  assign io_outputs_0_payload_0_pixel_10 = io_input_payload_0_pixel_10;
  assign io_outputs_0_payload_0_pixel_11 = io_input_payload_0_pixel_11;
  assign io_outputs_0_payload_0_pixel_12 = io_input_payload_0_pixel_12;
  assign io_outputs_0_payload_0_pixel_13 = io_input_payload_0_pixel_13;
  assign io_outputs_0_payload_0_pixel_14 = io_input_payload_0_pixel_14;
  assign io_outputs_0_payload_0_pixel_15 = io_input_payload_0_pixel_15;
  assign io_outputs_0_payload_0_endOfLine = io_input_payload_0_endOfLine;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && tmp_io_outputs_1_valid);
  assign io_outputs_1_payload_0_pixel_0 = io_input_payload_0_pixel_0;
  assign io_outputs_1_payload_0_pixel_1 = io_input_payload_0_pixel_1;
  assign io_outputs_1_payload_0_pixel_2 = io_input_payload_0_pixel_2;
  assign io_outputs_1_payload_0_pixel_3 = io_input_payload_0_pixel_3;
  assign io_outputs_1_payload_0_pixel_4 = io_input_payload_0_pixel_4;
  assign io_outputs_1_payload_0_pixel_5 = io_input_payload_0_pixel_5;
  assign io_outputs_1_payload_0_pixel_6 = io_input_payload_0_pixel_6;
  assign io_outputs_1_payload_0_pixel_7 = io_input_payload_0_pixel_7;
  assign io_outputs_1_payload_0_pixel_8 = io_input_payload_0_pixel_8;
  assign io_outputs_1_payload_0_pixel_9 = io_input_payload_0_pixel_9;
  assign io_outputs_1_payload_0_pixel_10 = io_input_payload_0_pixel_10;
  assign io_outputs_1_payload_0_pixel_11 = io_input_payload_0_pixel_11;
  assign io_outputs_1_payload_0_pixel_12 = io_input_payload_0_pixel_12;
  assign io_outputs_1_payload_0_pixel_13 = io_input_payload_0_pixel_13;
  assign io_outputs_1_payload_0_pixel_14 = io_input_payload_0_pixel_14;
  assign io_outputs_1_payload_0_pixel_15 = io_input_payload_0_pixel_15;
  assign io_outputs_1_payload_0_endOfLine = io_input_payload_0_endOfLine;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  always @(posedge clk) begin
    if(reset) begin
      tmp_io_outputs_0_valid <= 1'b1;
      tmp_io_outputs_1_valid <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        tmp_io_outputs_0_valid <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        tmp_io_outputs_1_valid <= 1'b0;
      end
      if(io_input_ready) begin
        tmp_io_outputs_0_valid <= 1'b1;
        tmp_io_outputs_1_valid <= 1'b1;
      end
    end
  end


endmodule

module StreamFork (
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_frame_line_pixel_0,
  input      [7:0]    io_input_payload_frame_line_pixel_1,
  input      [7:0]    io_input_payload_frame_line_pixel_2,
  input      [7:0]    io_input_payload_frame_line_pixel_3,
  input      [7:0]    io_input_payload_frame_line_pixel_4,
  input      [7:0]    io_input_payload_frame_line_pixel_5,
  input      [7:0]    io_input_payload_frame_line_pixel_6,
  input      [7:0]    io_input_payload_frame_line_pixel_7,
  input      [7:0]    io_input_payload_frame_line_pixel_8,
  input      [7:0]    io_input_payload_frame_line_pixel_9,
  input      [7:0]    io_input_payload_frame_line_pixel_10,
  input      [7:0]    io_input_payload_frame_line_pixel_11,
  input      [7:0]    io_input_payload_frame_line_pixel_12,
  input      [7:0]    io_input_payload_frame_line_pixel_13,
  input      [7:0]    io_input_payload_frame_line_pixel_14,
  input      [7:0]    io_input_payload_frame_line_pixel_15,
  input               io_input_payload_frame_line_endOfLine,
  input               io_input_payload_frame_endOfFrame,
  input               io_input_payload_endOfPack,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_0,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_1,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_2,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_3,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_4,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_5,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_6,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_7,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_8,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_9,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_10,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_11,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_12,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_13,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_14,
  output     [7:0]    io_outputs_0_payload_frame_line_pixel_15,
  output              io_outputs_0_payload_frame_line_endOfLine,
  output              io_outputs_0_payload_frame_endOfFrame,
  output              io_outputs_0_payload_endOfPack,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_0,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_1,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_2,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_3,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_4,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_5,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_6,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_7,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_8,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_9,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_10,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_11,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_12,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_13,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_14,
  output     [7:0]    io_outputs_1_payload_frame_line_pixel_15,
  output              io_outputs_1_payload_frame_line_endOfLine,
  output              io_outputs_1_payload_frame_endOfFrame,
  output              io_outputs_1_payload_endOfPack,
  input               clk,
  input               reset
);

  reg                 tmp_io_outputs_0_valid;
  reg                 tmp_io_outputs_1_valid;
  wire                when_Stream_l825;
  wire                when_Stream_l825_1;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l825) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l825_1) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l825 = ((! io_outputs_0_ready) && tmp_io_outputs_0_valid);
  assign when_Stream_l825_1 = ((! io_outputs_1_ready) && tmp_io_outputs_1_valid);
  assign io_outputs_0_valid = (io_input_valid && tmp_io_outputs_0_valid);
  assign io_outputs_0_payload_frame_line_pixel_0 = io_input_payload_frame_line_pixel_0;
  assign io_outputs_0_payload_frame_line_pixel_1 = io_input_payload_frame_line_pixel_1;
  assign io_outputs_0_payload_frame_line_pixel_2 = io_input_payload_frame_line_pixel_2;
  assign io_outputs_0_payload_frame_line_pixel_3 = io_input_payload_frame_line_pixel_3;
  assign io_outputs_0_payload_frame_line_pixel_4 = io_input_payload_frame_line_pixel_4;
  assign io_outputs_0_payload_frame_line_pixel_5 = io_input_payload_frame_line_pixel_5;
  assign io_outputs_0_payload_frame_line_pixel_6 = io_input_payload_frame_line_pixel_6;
  assign io_outputs_0_payload_frame_line_pixel_7 = io_input_payload_frame_line_pixel_7;
  assign io_outputs_0_payload_frame_line_pixel_8 = io_input_payload_frame_line_pixel_8;
  assign io_outputs_0_payload_frame_line_pixel_9 = io_input_payload_frame_line_pixel_9;
  assign io_outputs_0_payload_frame_line_pixel_10 = io_input_payload_frame_line_pixel_10;
  assign io_outputs_0_payload_frame_line_pixel_11 = io_input_payload_frame_line_pixel_11;
  assign io_outputs_0_payload_frame_line_pixel_12 = io_input_payload_frame_line_pixel_12;
  assign io_outputs_0_payload_frame_line_pixel_13 = io_input_payload_frame_line_pixel_13;
  assign io_outputs_0_payload_frame_line_pixel_14 = io_input_payload_frame_line_pixel_14;
  assign io_outputs_0_payload_frame_line_pixel_15 = io_input_payload_frame_line_pixel_15;
  assign io_outputs_0_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_0_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_0_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && tmp_io_outputs_1_valid);
  assign io_outputs_1_payload_frame_line_pixel_0 = io_input_payload_frame_line_pixel_0;
  assign io_outputs_1_payload_frame_line_pixel_1 = io_input_payload_frame_line_pixel_1;
  assign io_outputs_1_payload_frame_line_pixel_2 = io_input_payload_frame_line_pixel_2;
  assign io_outputs_1_payload_frame_line_pixel_3 = io_input_payload_frame_line_pixel_3;
  assign io_outputs_1_payload_frame_line_pixel_4 = io_input_payload_frame_line_pixel_4;
  assign io_outputs_1_payload_frame_line_pixel_5 = io_input_payload_frame_line_pixel_5;
  assign io_outputs_1_payload_frame_line_pixel_6 = io_input_payload_frame_line_pixel_6;
  assign io_outputs_1_payload_frame_line_pixel_7 = io_input_payload_frame_line_pixel_7;
  assign io_outputs_1_payload_frame_line_pixel_8 = io_input_payload_frame_line_pixel_8;
  assign io_outputs_1_payload_frame_line_pixel_9 = io_input_payload_frame_line_pixel_9;
  assign io_outputs_1_payload_frame_line_pixel_10 = io_input_payload_frame_line_pixel_10;
  assign io_outputs_1_payload_frame_line_pixel_11 = io_input_payload_frame_line_pixel_11;
  assign io_outputs_1_payload_frame_line_pixel_12 = io_input_payload_frame_line_pixel_12;
  assign io_outputs_1_payload_frame_line_pixel_13 = io_input_payload_frame_line_pixel_13;
  assign io_outputs_1_payload_frame_line_pixel_14 = io_input_payload_frame_line_pixel_14;
  assign io_outputs_1_payload_frame_line_pixel_15 = io_input_payload_frame_line_pixel_15;
  assign io_outputs_1_payload_frame_line_endOfLine = io_input_payload_frame_line_endOfLine;
  assign io_outputs_1_payload_frame_endOfFrame = io_input_payload_frame_endOfFrame;
  assign io_outputs_1_payload_endOfPack = io_input_payload_endOfPack;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  always @(posedge clk) begin
    if(reset) begin
      tmp_io_outputs_0_valid <= 1'b1;
      tmp_io_outputs_1_valid <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        tmp_io_outputs_0_valid <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        tmp_io_outputs_1_valid <= 1'b0;
      end
      if(io_input_ready) begin
        tmp_io_outputs_0_valid <= 1'b1;
        tmp_io_outputs_1_valid <= 1'b1;
      end
    end
  end


endmodule

module StreamFifoHighPerf (
  input               push_valid,
  output              push_ready,
  input      [7:0]    push_payload_0_pixel_0,
  input      [7:0]    push_payload_0_pixel_1,
  input      [7:0]    push_payload_0_pixel_2,
  input      [7:0]    push_payload_0_pixel_3,
  input      [7:0]    push_payload_0_pixel_4,
  input      [7:0]    push_payload_0_pixel_5,
  input      [7:0]    push_payload_0_pixel_6,
  input      [7:0]    push_payload_0_pixel_7,
  input      [7:0]    push_payload_0_pixel_8,
  input      [7:0]    push_payload_0_pixel_9,
  input      [7:0]    push_payload_0_pixel_10,
  input      [7:0]    push_payload_0_pixel_11,
  input      [7:0]    push_payload_0_pixel_12,
  input      [7:0]    push_payload_0_pixel_13,
  input      [7:0]    push_payload_0_pixel_14,
  input      [7:0]    push_payload_0_pixel_15,
  input               push_payload_0_endOfLine,
  output              pop_valid,
  input               pop_ready,
  output     [7:0]    pop_payload_0_pixel_0,
  output     [7:0]    pop_payload_0_pixel_1,
  output     [7:0]    pop_payload_0_pixel_2,
  output     [7:0]    pop_payload_0_pixel_3,
  output     [7:0]    pop_payload_0_pixel_4,
  output     [7:0]    pop_payload_0_pixel_5,
  output     [7:0]    pop_payload_0_pixel_6,
  output     [7:0]    pop_payload_0_pixel_7,
  output     [7:0]    pop_payload_0_pixel_8,
  output     [7:0]    pop_payload_0_pixel_9,
  output     [7:0]    pop_payload_0_pixel_10,
  output     [7:0]    pop_payload_0_pixel_11,
  output     [7:0]    pop_payload_0_pixel_12,
  output     [7:0]    pop_payload_0_pixel_13,
  output     [7:0]    pop_payload_0_pixel_14,
  output     [7:0]    pop_payload_0_pixel_15,
  output              pop_payload_0_endOfLine,
  input               flush,
  input               clk,
  input               reset
);

  reg        [128:0]  tmp_ram_port0;
  wire       [8:0]    tmp_pushPtr_valueNext;
  wire       [0:0]    tmp_pushPtr_valueNext_1;
  wire       [8:0]    tmp_popPtr_valueNext;
  wire       [0:0]    tmp_popPtr_valueNext_1;
  wire       [128:0]  tmp_ram_port;
  reg                 tmp_1;
  wire                popEvent_valid;
  reg                 popEvent_ready;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [8:0]    pushPtr_valueNext;
  reg        [8:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [8:0]    popPtr_valueNext;
  reg        [8:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                pushing;
  wire                popping;
  wire                empty;
  wire                full;
  reg                 tmp_popEvent_valid;
  reg                 rValid;
  wire       [7:0]    rData_0_pixel_0;
  wire       [7:0]    rData_0_pixel_1;
  wire       [7:0]    rData_0_pixel_2;
  wire       [7:0]    rData_0_pixel_3;
  wire       [7:0]    rData_0_pixel_4;
  wire       [7:0]    rData_0_pixel_5;
  wire       [7:0]    rData_0_pixel_6;
  wire       [7:0]    rData_0_pixel_7;
  wire       [7:0]    rData_0_pixel_8;
  wire       [7:0]    rData_0_pixel_9;
  wire       [7:0]    rData_0_pixel_10;
  wire       [7:0]    rData_0_pixel_11;
  wire       [7:0]    rData_0_pixel_12;
  wire       [7:0]    rData_0_pixel_13;
  wire       [7:0]    rData_0_pixel_14;
  wire       [7:0]    rData_0_pixel_15;
  wire                rData_0_endOfLine;
  wire       [128:0]  tmp_rData_0_pixel_0;
  wire       [127:0]  tmp_rData_0_pixel_0_1;
  wire                when_StreamFifoHighPerf_l38;
  wire                when_StreamFifoHighPerf_l42;
  reg [128:0] ram [0:511];

  assign tmp_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign tmp_pushPtr_valueNext = {8'd0, tmp_pushPtr_valueNext_1};
  assign tmp_popPtr_valueNext_1 = popPtr_willIncrement;
  assign tmp_popPtr_valueNext = {8'd0, tmp_popPtr_valueNext_1};
  assign tmp_ram_port = {push_payload_0_endOfLine,{push_payload_0_pixel_15,{push_payload_0_pixel_14,{push_payload_0_pixel_13,{push_payload_0_pixel_12,{push_payload_0_pixel_11,{push_payload_0_pixel_10,{push_payload_0_pixel_9,{push_payload_0_pixel_8,{push_payload_0_pixel_7,{push_payload_0_pixel_6,{push_payload_0_pixel_5,{push_payload_0_pixel_4,{push_payload_0_pixel_3,{push_payload_0_pixel_2,{push_payload_0_pixel_1,push_payload_0_pixel_0}}}}}}}}}}}}}}}};
  always @(posedge clk) begin
    if(popEvent_ready) begin
      tmp_ram_port0 <= ram[popPtr_value];
    end
  end

  always @(posedge clk) begin
    if(tmp_1) begin
      ram[pushPtr_value] <= tmp_ram_port;
    end
  end

  always @(*) begin
    tmp_1 = 1'b0;
    if(pushing) begin
      tmp_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 9'h1ff);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + tmp_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 9'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 9'h1ff);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + tmp_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 9'h0;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign pushing = (push_valid && push_ready);
  assign popping = (popEvent_valid && popEvent_ready);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign push_ready = (! full);
  assign popEvent_valid = ((! empty) && (! (tmp_popEvent_valid && (! full))));
  assign tmp_rData_0_pixel_0 = tmp_ram_port0[128 : 0];
  assign tmp_rData_0_pixel_0_1 = tmp_rData_0_pixel_0[127 : 0];
  assign rData_0_pixel_0 = tmp_rData_0_pixel_0_1[7 : 0];
  assign rData_0_pixel_1 = tmp_rData_0_pixel_0_1[15 : 8];
  assign rData_0_pixel_2 = tmp_rData_0_pixel_0_1[23 : 16];
  assign rData_0_pixel_3 = tmp_rData_0_pixel_0_1[31 : 24];
  assign rData_0_pixel_4 = tmp_rData_0_pixel_0_1[39 : 32];
  assign rData_0_pixel_5 = tmp_rData_0_pixel_0_1[47 : 40];
  assign rData_0_pixel_6 = tmp_rData_0_pixel_0_1[55 : 48];
  assign rData_0_pixel_7 = tmp_rData_0_pixel_0_1[63 : 56];
  assign rData_0_pixel_8 = tmp_rData_0_pixel_0_1[71 : 64];
  assign rData_0_pixel_9 = tmp_rData_0_pixel_0_1[79 : 72];
  assign rData_0_pixel_10 = tmp_rData_0_pixel_0_1[87 : 80];
  assign rData_0_pixel_11 = tmp_rData_0_pixel_0_1[95 : 88];
  assign rData_0_pixel_12 = tmp_rData_0_pixel_0_1[103 : 96];
  assign rData_0_pixel_13 = tmp_rData_0_pixel_0_1[111 : 104];
  assign rData_0_pixel_14 = tmp_rData_0_pixel_0_1[119 : 112];
  assign rData_0_pixel_15 = tmp_rData_0_pixel_0_1[127 : 120];
  assign rData_0_endOfLine = tmp_rData_0_pixel_0[128];
  always @(*) begin
    popEvent_ready = pop_ready;
    if(when_StreamFifoHighPerf_l38) begin
      popEvent_ready = 1'b1;
    end
  end

  assign when_StreamFifoHighPerf_l38 = (! rValid);
  assign pop_valid = rValid;
  assign pop_payload_0_pixel_0 = rData_0_pixel_0;
  assign pop_payload_0_pixel_1 = rData_0_pixel_1;
  assign pop_payload_0_pixel_2 = rData_0_pixel_2;
  assign pop_payload_0_pixel_3 = rData_0_pixel_3;
  assign pop_payload_0_pixel_4 = rData_0_pixel_4;
  assign pop_payload_0_pixel_5 = rData_0_pixel_5;
  assign pop_payload_0_pixel_6 = rData_0_pixel_6;
  assign pop_payload_0_pixel_7 = rData_0_pixel_7;
  assign pop_payload_0_pixel_8 = rData_0_pixel_8;
  assign pop_payload_0_pixel_9 = rData_0_pixel_9;
  assign pop_payload_0_pixel_10 = rData_0_pixel_10;
  assign pop_payload_0_pixel_11 = rData_0_pixel_11;
  assign pop_payload_0_pixel_12 = rData_0_pixel_12;
  assign pop_payload_0_pixel_13 = rData_0_pixel_13;
  assign pop_payload_0_pixel_14 = rData_0_pixel_14;
  assign pop_payload_0_pixel_15 = rData_0_pixel_15;
  assign pop_payload_0_endOfLine = rData_0_endOfLine;
  assign when_StreamFifoHighPerf_l42 = (pushing != popping);
  always @(posedge clk) begin
    if(reset) begin
      pushPtr_value <= 9'h0;
      popPtr_value <= 9'h0;
      risingOccupancy <= 1'b0;
      tmp_popEvent_valid <= 1'b0;
      rValid <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      tmp_popEvent_valid <= (popPtr_valueNext == pushPtr_value);
      if(popEvent_ready) begin
        rValid <= popEvent_valid;
      end
      if(when_StreamFifoHighPerf_l42) begin
        risingOccupancy <= pushing;
      end
      if(flush) begin
        rValid <= 1'b0;
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
